

module sa_acc
(
  input clk,
  input rst,
  input start,
  input [1-1:0] acc_user_done_rd_data,
  input [1-1:0] acc_user_done_wr_data,
  output [1-1:0] acc_user_request_read,
  input [1-1:0] acc_user_read_data_valid,
  input [32-1:0] acc_user_read_data,
  input [1-1:0] acc_user_available_write,
  output [1-1:0] acc_user_request_write,
  output [32-1:0] acc_user_write_data,
  output acc_user_done
);

  reg start_reg;
  wire [1-1:0] sa_aws_done;
  assign acc_user_done = &sa_aws_done;

  always @(posedge clk) begin
    if(rst) begin
      start_reg <= 0;
    end else begin
      start_reg <= start_reg | start;
    end
  end

  (* keep_hierarchy = "yes" *)

  sa_aws
  sa_aws_0
  (
    .clk(clk),
    .rst(rst),
    .start(start_reg),
    .sa_aws_done_rd_data(acc_user_done_rd_data[0]),
    .sa_aws_done_wr_data(acc_user_done_wr_data[0]),
    .sa_aws_request_read(acc_user_request_read[0]),
    .sa_aws_read_data_valid(acc_user_read_data_valid[0]),
    .sa_aws_read_data(acc_user_read_data[31:0]),
    .sa_aws_available_write(acc_user_available_write[0]),
    .sa_aws_request_write(acc_user_request_write[0]),
    .sa_aws_write_data(acc_user_write_data[31:0]),
    .sa_aws_done(sa_aws_done[0])
  );


  initial begin
    start_reg = 0;
  end


endmodule



module sa_aws
(
  input clk,
  input rst,
  input start,
  input sa_aws_done_rd_data,
  input sa_aws_done_wr_data,
  output sa_aws_request_read,
  input sa_aws_read_data_valid,
  input [32-1:0] sa_aws_read_data,
  input sa_aws_available_write,
  output reg sa_aws_request_write,
  output reg [32-1:0] sa_aws_write_data,
  output sa_aws_done
);

  assign sa_aws_done = &{ sa_aws_done_wr_data, sa_aws_done_rd_data };
  reg start_pipe;
  reg pop_data;
  wire available_pop;
  wire [16-1:0] data_out;
  reg [16-1:0] config_data;
  reg [2-1:0] fms_sd;
  localparam [2-1:0] fsm_sd_idle = 0;
  localparam [2-1:0] fsm_sd_send_data = 1;
  localparam [2-1:0] fsm_sd_done = 2;
  reg flag;
  wire sa_done;
  reg sa_rd;
  reg [10-1:0] sa_rd_addr;
  wire sa_out_v;
  wire [7-1:0] sa_out_data;

  always @(posedge clk) begin
    if(rst) begin
      pop_data <= 0;
      fms_sd <= fsm_sd_idle;
      flag <= 0;
    end else begin
      if(start) begin
        start_pipe <= 0;
        pop_data <= 0;
        flag <= 0;
        case(fms_sd)
          fsm_sd_idle: begin
            if(available_pop) begin
              pop_data <= 1;
              flag <= 1;
              fms_sd <= fsm_sd_send_data;
            end 
          end
          fsm_sd_send_data: begin
            config_data <= data_out;
            fms_sd <= fsm_sd_done;
          end
          fsm_sd_done: begin
            start_pipe <= 1;
          end
        endcase
      end 
    end
  end


  //Data Consumer - Begin
  reg [2-1:0] fsm_consume;
  localparam fsm_consume_wait = 0;
  localparam fsm_consume_consume = 1;
  localparam fsm_consume_verify = 2;
  localparam fsm_consume_done = 3;

  always @(posedge clk) begin
    if(rst) begin
      sa_rd <= 0;
      sa_rd_addr <= 0;
      sa_aws_request_write <= 0;
      fsm_consume <= fsm_consume_wait;
    end else begin
      sa_rd <= 0;
      sa_aws_request_write <= 0;
      case(fsm_consume)
        fsm_consume_wait: begin
          if(sa_aws_available_write) begin
            if(sa_done) begin
              sa_rd <= 1;
              fsm_consume <= fsm_consume_consume;
            end 
          end 
        end
        fsm_consume_consume: begin
          if(sa_out_v) begin
            sa_aws_request_write <= 1;
            sa_aws_write_data <= { 25'd0, sa_out_data };
            sa_rd_addr <= sa_rd_addr + 1;
            fsm_consume <= fsm_consume_verify;
          end 
        end
        fsm_consume_verify: begin
          if(sa_rd_addr == 512) begin
            fsm_consume <= fsm_consume_done;
          end else begin
            fsm_consume <= fsm_consume_wait;
          end
        end
        fsm_consume_done: begin
        end
      endcase
    end
  end

  //Data Consumer - Begin
  (* keep_hierarchy = "yes" *)

  fecth_data_32_16
  fecth_data_32_16
  (
    .clk(clk),
    .rst(rst),
    .start(start),
    .request_read(sa_aws_request_read),
    .data_valid(sa_aws_read_data_valid),
    .read_data(sa_aws_read_data),
    .pop_data(pop_data),
    .available_pop(available_pop),
    .data_out(data_out)
  );


  sa_pipeline_6th_64cells
  sa_pipeline_6th_64cells
  (
    .clk(clk),
    .rst(rst),
    .start(start_pipe),
    .n_exec(config_data),
    .done(sa_done),
    .rd(sa_rd),
    .rd_addr(sa_rd_addr[8:0]),
    .out_v(sa_out_v),
    .out_data(sa_out_data)
  );


  initial begin
    sa_aws_request_write = 0;
    sa_aws_write_data = 0;
    start_pipe = 0;
    pop_data = 0;
    config_data = 0;
    fms_sd = 0;
    flag = 0;
    sa_rd = 0;
    sa_rd_addr = 0;
    fsm_consume = 0;
  end


endmodule



module fecth_data_32_16
(
  input clk,
  input start,
  input rst,
  output reg request_read,
  input data_valid,
  input [32-1:0] read_data,
  input pop_data,
  output reg available_pop,
  output [16-1:0] data_out
);

  reg [1-1:0] fsm_read;
  reg [1-1:0] fsm_control;
  reg [32-1:0] data;
  reg [32-1:0] buffer;
  reg [2-1:0] count;
  reg has_buffer;
  reg buffer_read;
  reg en;

  assign data_out = data[15:0];

  always @(posedge clk) begin
    if(rst) begin
      en <= 1'b0;
    end else begin
      en <= (en)? en : start;
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      fsm_read <= 0;
      request_read <= 0;
      has_buffer <= 0;
    end else begin
      request_read <= 0;
      case(fsm_read)
        0: begin
          if(en & data_valid) begin
            buffer <= read_data;
            request_read <= 1;
            has_buffer <= 1;
            fsm_read <= 1;
          end 
        end
        1: begin
          if(buffer_read) begin
            has_buffer <= 0;
            fsm_read <= 0;
          end 
        end
      endcase
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      fsm_control <= 0;
      available_pop <= 0;
      count <= 0;
      buffer_read <= 0;
    end else begin
      buffer_read <= 0;
      case(fsm_control)
        0: begin
          if(has_buffer) begin
            data <= buffer;
            count <= 1;
            buffer_read <= 1;
            available_pop <= 1;
            fsm_control <= 1;
          end 
        end
        1: begin
          if(pop_data & ~count[1]) begin
            count <= count << 1;
            data <= data[31:16];
          end 
          if(pop_data & count[1] & has_buffer) begin
            count <= 1;
            data <= buffer;
            buffer_read <= 1;
          end 
          if(count[1] & pop_data & ~has_buffer) begin
            count <= count << 1;
            data <= data[31:16];
            available_pop <= 0;
            fsm_control <= 0;
          end 
        end
      endcase
    end
  end


  initial begin
    request_read = 0;
    available_pop = 0;
    fsm_read = 0;
    fsm_control = 0;
    data = 0;
    buffer = 0;
    count = 0;
    has_buffer = 0;
    buffer_read = 0;
    en = 0;
  end


endmodule



module sa_pipeline_6th_64cells
(
  input clk,
  input rst,
  input start,
  input [16-1:0] n_exec,
  output reg done,
  input rd,
  input [9-1:0] rd_addr,
  output out_v,
  output [7-1:0] out_data
);

  // basic control inputs
  // -----
  wire pipe_start;
  reg [17-1:0] counter_total;
  // Threads controller output wires
  wire [3-1:0] th_idx;
  wire th_v;
  wire [6-1:0] th_ca;
  wire [6-1:0] th_cb;
  // -----

  always @(posedge clk) begin
    if(rst) begin
      counter_total <= 0;
      done <= 0;
    end else begin
      if(pipe_start) begin
        if((th_idx == 5) && ~th_v && &{ th_ca, th_cb }) begin
          counter_total <= counter_total + 1;
        end 
        if(counter_total == n_exec) begin
          done <= 1;
        end 
      end 
    end
  end

  // st1 output wires
  wire st1_rdy;
  wire [3-1:0] st1_idx;
  wire st1_v;
  wire [6-1:0] st1_ca;
  wire [6-1:0] st1_cb;
  wire [6-1:0] st1_na;
  wire st1_na_v;
  wire [6-1:0] st1_nb;
  wire st1_nb_v;
  wire st1_sw;
  wire [16-1:0] st1_wa;
  wire [16-1:0] st1_wb;
  // -----
  // st2 output wires
  wire [3-1:0] st2_idx;
  wire st2_v;
  wire [6-1:0] st2_ca;
  wire [6-1:0] st2_cb;
  wire [6-1:0] st2_na;
  wire st2_na_v;
  wire [6-1:0] st2_nb;
  wire st2_nb_v;
  wire [24-1:0] st2_va;
  wire [4-1:0] st2_va_v;
  wire [24-1:0] st2_vb;
  wire [4-1:0] st2_vb_v;
  wire st2_sw;
  wire [16-1:0] st2_wa;
  wire [16-1:0] st2_wb;
  // -----
  // st3 output wires
  wire [3-1:0] st3_idx;
  wire st3_v;
  wire [6-1:0] st3_ca;
  wire [6-1:0] st3_cb;
  wire [24-1:0] st3_cva;
  wire [4-1:0] st3_cva_v;
  wire [24-1:0] st3_cvb;
  wire [4-1:0] st3_cvb_v;
  wire [16-1:0] st3_wb;
  // -----
  // st4 output wires
  wire [3-1:0] st4_idx;
  wire st4_v;
  wire [6-1:0] st4_ca;
  wire [6-1:0] st4_cb;
  wire [24-1:0] st4_cva;
  wire [4-1:0] st4_cva_v;
  wire [24-1:0] st4_cvb;
  wire [4-1:0] st4_cvb_v;
  wire [36-1:0] st4_dvac;
  wire [36-1:0] st4_dvbc;
  // -----
  // st5 output wires
  wire [3-1:0] st5_idx;
  wire st5_v;
  wire [18-1:0] st5_dvac;
  wire [18-1:0] st5_dvbc;
  wire [36-1:0] st5_dvas;
  wire [36-1:0] st5_dvbs;
  // -----
  // st6 output wires
  wire [3-1:0] st6_idx;
  wire st6_v;
  wire [9-1:0] st6_dvac;
  wire [9-1:0] st6_dvbc;
  wire [18-1:0] st6_dvas;
  wire [18-1:0] st6_dvbs;
  // -----
  // st7 output wires
  wire [3-1:0] st7_idx;
  wire st7_v;
  wire [9-1:0] st7_dc;
  wire [9-1:0] st7_dvas;
  wire [9-1:0] st7_dvbs;
  // st8 output wires
  wire [3-1:0] st8_idx;
  wire st8_v;
  wire [9-1:0] st8_dc;
  wire [9-1:0] st8_ds;
  // -----
  // st9 output wires
  wire [3-1:0] st9_idx;
  wire st9_v;
  wire st9_sw;
  // -----
  // st10 output wires
  wire [3-1:0] st10_idx;
  wire st10_v;
  wire st10_sw;
  // -----
  assign pipe_start = &{ start, st1_rdy };

  th_controller_6th_64cells
  th_controller_6th_64cells
  (
    .clk(clk),
    .rst(rst),
    .start(pipe_start),
    .done(done),
    .idx_out(th_idx),
    .v_out(th_v),
    .ca_out(th_ca),
    .cb_out(th_cb)
  );


  st1_c2n_6th_64cells
  st1_c2n_6th_64cells
  (
    .rd(rd),
    .rd_addr(rd_addr),
    .out_v(out_v),
    .out_data(out_data),
    .clk(clk),
    .rst(rst),
    .rdy(st1_rdy),
    .idx_in(th_idx),
    .v_in(th_v),
    .ca_in(th_ca),
    .cb_in(th_cb),
    .sw_in(st10_sw),
    .st1_wb_in(st1_wb),
    .idx_out(st1_idx),
    .v_out(st1_v),
    .ca_out(st1_ca),
    .cb_out(st1_cb),
    .na_out(st1_na),
    .na_v_out(st1_na_v),
    .nb_out(st1_nb),
    .nb_v_out(st1_nb_v),
    .sw_out(st1_sw),
    .wa_out(st1_wa),
    .wb_out(st1_wb)
  );


  st2_n_6th_64cells
  st2_n_6th_64cells
  (
    .clk(clk),
    .idx_in(st1_idx),
    .v_in(st1_v),
    .ca_in(st1_ca),
    .cb_in(st1_cb),
    .na_in(st1_na),
    .na_v_in(st1_na_v),
    .nb_in(st1_nb),
    .nb_v_in(st1_nb_v),
    .sw_in(st1_sw),
    .wa_in(st1_wa),
    .wb_in(st1_wb),
    .idx_out(st2_idx),
    .v_out(st2_v),
    .ca_out(st2_ca),
    .cb_out(st2_cb),
    .na_out(st2_na),
    .na_v_out(st2_na_v),
    .nb_out(st2_nb),
    .nb_v_out(st2_nb_v),
    .va_out(st2_va),
    .va_v_out(st2_va_v),
    .vb_out(st2_vb),
    .vb_v_out(st2_vb_v),
    .sw_out(st2_sw),
    .wa_out(st2_wa),
    .wb_out(st2_wb)
  );


  st3_n2c_6th_64cells
  st3_n2c_6th_64cells
  (
    .clk(clk),
    .rst(rst),
    .idx_in(st2_idx),
    .v_in(st2_v),
    .ca_in(st2_ca),
    .cb_in(st2_cb),
    .na_in(st2_na),
    .na_v_in(st2_na_v),
    .nb_in(st2_nb),
    .nb_v_in(st2_nb_v),
    .va_in(st2_va),
    .va_v_in(st2_va_v),
    .vb_in(st2_vb),
    .vb_v_in(st2_vb_v),
    .st3_wb_in(st3_wb),
    .sw_in(st2_sw),
    .wa_in(st2_wa),
    .wb_in(st2_wb),
    .idx_out(st3_idx),
    .v_out(st3_v),
    .ca_out(st3_ca),
    .cb_out(st3_cb),
    .cva_out(st3_cva),
    .cva_v_out(st3_cva_v),
    .cvb_out(st3_cvb),
    .cvb_v_out(st3_cvb_v),
    .wb_out(st3_wb)
  );


  st4_d1_6th_64cells
  st4_d1_6th_64cells
  (
    .clk(clk),
    .idx_in(st3_idx),
    .v_in(st3_v),
    .ca_in(st3_ca),
    .cb_in(st3_cb),
    .cva_in(st3_cva),
    .cva_v_in(st3_cva_v),
    .cvb_in(st3_cvb),
    .cvb_v_in(st3_cvb_v),
    .idx_out(st4_idx),
    .v_out(st4_v),
    .ca_out(st4_ca),
    .cb_out(st4_cb),
    .cva_out(st4_cva),
    .cva_v_out(st4_cva_v),
    .cvb_out(st4_cvb),
    .cvb_v_out(st4_cvb_v),
    .dvac_out(st4_dvac),
    .dvbc_out(st4_dvbc)
  );


  st5_d2_s1_6th_64cells
  st5_d2_s1_6th_64cells
  (
    .clk(clk),
    .idx_in(st4_idx),
    .v_in(st4_v),
    .ca_in(st4_ca),
    .cb_in(st4_cb),
    .cva_in(st4_cva),
    .cva_v_in(st4_cva_v),
    .cvb_in(st4_cvb),
    .cvb_v_in(st4_cvb_v),
    .dvac_in(st4_dvac),
    .dvbc_in(st4_dvbc),
    .idx_out(st5_idx),
    .v_out(st5_v),
    .dvac_out(st5_dvac),
    .dvbc_out(st5_dvbc),
    .dvas_out(st5_dvas),
    .dvbs_out(st5_dvbs)
  );


  st6_s2_6th_64cells
  st6_s2_6th_64cells
  (
    .clk(clk),
    .idx_in(st5_idx),
    .v_in(st5_v),
    .dvac_in(st5_dvac),
    .dvbc_in(st5_dvbc),
    .dvas_in(st5_dvas),
    .dvbs_in(st5_dvbs),
    .idx_out(st6_idx),
    .v_out(st6_v),
    .dvac_out(st6_dvac),
    .dvbc_out(st6_dvbc),
    .dvas_out(st6_dvas),
    .dvbs_out(st6_dvbs)
  );


  st7_s3_6th_64cells
  st7_s3_6th_64cells
  (
    .clk(clk),
    .idx_in(st6_idx),
    .v_in(st6_v),
    .dvac_in(st6_dvac),
    .dvbc_in(st6_dvbc),
    .dvas_in(st6_dvas),
    .dvbs_in(st6_dvbs),
    .idx_out(st7_idx),
    .v_out(st7_v),
    .dc_out(st7_dc),
    .dvas_out(st7_dvas),
    .dvbs_out(st7_dvbs)
  );


  st8_s4_6th_64cells
  st8_s4_6th_64cells
  (
    .clk(clk),
    .idx_in(st7_idx),
    .v_in(st7_v),
    .dc_in(st7_dc),
    .dvas_in(st7_dvas),
    .dvbs_in(st7_dvbs),
    .idx_out(st8_idx),
    .v_out(st8_v),
    .dc_out(st8_dc),
    .ds_out(st8_ds)
  );


  st9_cmp_6th_64cells
  st9_cmp_6th_64cells
  (
    .clk(clk),
    .idx_in(st8_idx),
    .v_in(st8_v),
    .dc_in(st8_dc),
    .ds_in(st8_ds),
    .idx_out(st9_idx),
    .v_out(st9_v),
    .sw_out(st9_sw)
  );


  st10_reg_6th_64cells
  st10_reg_6th_64cells
  (
    .clk(clk),
    .idx_in(st9_idx),
    .v_in(st9_v),
    .sw_in(st9_sw),
    .idx_out(st10_idx),
    .v_out(st10_v),
    .sw_out(st10_sw)
  );


  initial begin
    done = 0;
    counter_total = 0;
  end


endmodule



module th_controller_6th_64cells
(
  input clk,
  input rst,
  input start,
  input done,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [6-1:0] ca_out,
  output reg [6-1:0] cb_out
);

  reg [6-1:0] flag_f_exec;
  reg [6-1:0] v_r;
  reg [3-1:0] idx_r;
  wire [12-1:0] counter;
  wire [12-1:0] counter_t;
  wire [12-1:0] counter_wr;
  wire [6-1:0] ca_out_t;
  wire [6-1:0] cb_out_t;
  assign counter_t = (flag_f_exec[idx_r])? 0 : counter;
  assign counter_wr = (&counter_t)? 0 : counter_t + 1;
  assign ca_out_t = counter_t[5:0];
  assign cb_out_t = counter_t[11:6];

  always @(posedge clk) begin
    if(rst) begin
      idx_out <= 0;
      v_out <= 0;
      ca_out <= 0;
      cb_out <= 0;
      idx_r <= 0;
      flag_f_exec <= 6'b111111;
      v_r <= 6'b111111;
    end else begin
      if(start) begin
        idx_out <= idx_r;
        v_out <= (done)? 1'b0 : v_r[idx_r];
        ca_out <= ca_out_t;
        cb_out <= cb_out_t;
        v_r[idx_r] <= ~v_r[idx_r];
        if(!v_r[idx_r]) begin
          flag_f_exec[idx_r] <= 0;
          if(idx_r == 5) begin
            idx_r <= 0;
          end else begin
            idx_r <= idx_r + 1;
          end
        end 
      end 
    end
  end


  mem_2r_1w_width12_depth3
  #(
    .init_file("./th.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width12_depth3
  (
    .clk(clk),
    .rd_addr0(idx_r),
    .out0(counter),
    .wr(~v_r[idx_r]),
    .wr_addr(idx_r),
    .wr_data(counter_wr)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    flag_f_exec = 0;
    v_r = 0;
    idx_r = 0;
  end


endmodule



module mem_2r_1w_width12_depth3 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [3-1:0] rd_addr0,
  input [3-1:0] rd_addr1,
  output [12-1:0] out0,
  output [12-1:0] out1,
  input wr,
  input [3-1:0] wr_addr,
  input [12-1:0] wr_data
);

  (*rom_style = "block" *) reg [12-1:0] mem[0:2**3-1];
  /*
  reg [12-1:0] mem [0:2**3-1];
  */
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end

  //synthesis translate_on

  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end


endmodule



module st1_c2n_6th_64cells
(
  input clk,
  input rst,
  input rd,
  input [9-1:0] rd_addr,
  output reg out_v,
  output reg [7-1:0] out_data,
  input [3-1:0] idx_in,
  input v_in,
  input [6-1:0] ca_in,
  input [6-1:0] cb_in,
  input sw_in,
  input [16-1:0] st1_wb_in,
  output reg rdy,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [6-1:0] ca_out,
  output reg [6-1:0] cb_out,
  output reg [6-1:0] na_out,
  output reg na_v_out,
  output reg [6-1:0] nb_out,
  output reg nb_v_out,
  output reg sw_out,
  output reg [16-1:0] wa_out,
  output reg [16-1:0] wb_out
);

  reg flag;
  reg [4-1:0] counter;
  reg fifo_init;
  wire [6-1:0] na_t;
  wire na_v_t;
  wire [6-1:0] nb_t;
  wire nb_v_t;
  wire [16-1:0] wa_t;
  wire [16-1:0] wb_t;
  wire fifoa_wr_en;
  wire fifoa_rd_en;
  wire [16-1:0] fifoa_data;
  wire fifob_wr_en;
  wire fifob_rd_en;
  wire [16-1:0] fifob_data;
  wire [3-1:0] wa_idx;
  wire [6-1:0] wa_c;
  wire [6-1:0] wa_n;
  wire wa_n_v;
  wire [3-1:0] wb_idx;
  wire [6-1:0] wb_c;
  wire [6-1:0] wb_n;
  wire wb_n_v;
  wire m_wr;
  wire [9-1:0] m_wr_addr;
  wire [7-1:0] m_wr_data;
  assign fifoa_data = { idx_in, ca_in, nb_v_t, nb_t };
  assign fifob_data = { idx_in, cb_in, na_v_t, na_t };
  assign fifoa_rd_en = &{ rdy, v_in };
  assign fifob_rd_en = &{ rdy, v_in };
  assign fifoa_wr_en = |{ &{ rdy, v_in }, fifo_init };
  assign fifob_wr_en = |{ &{ rdy, v_in }, fifo_init };
  assign wa_n = wa_t[5:0];
  assign wa_n_v = wa_t[6];
  assign wa_c = wa_t[12:7];
  assign wa_idx = wa_t[15:13];
  assign wb_n = st1_wb_in[5:0];
  assign wb_n_v = st1_wb_in[6];
  assign wb_c = st1_wb_in[12:7];
  assign wb_idx = st1_wb_in[15:13];
  assign m_wr = sw_in;
  assign m_wr_addr = (flag)? { wa_idx, wa_c } : { wb_idx, wb_c };
  assign m_wr_data = (flag)? { wa_n_v, wa_n } : { wb_n_v, wb_n };

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    na_out <= na_t;
    na_v_out <= na_v_t;
    nb_out <= nb_t;
    nb_v_out <= nb_v_t;
    sw_out <= sw_in;
    wa_out <= wa_t;
    wb_out <= wb_t;
    out_v <= rd;
    out_data <= { na_v_t, na_t };
  end


  always @(posedge clk) begin
    if(rst) begin
      flag <= 1;
    end else begin
      if(sw_in) begin
        flag <= ~flag;
      end 
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      rdy <= 0;
      fifo_init <= 0;
      counter <= 0;
    end else begin
      if(counter == 4) begin
        rdy <= 1;
        fifo_init <= 0;
      end else begin
        counter <= counter + 1;
        fifo_init <= 1;
      end
    end
  end


  mem_2r_1w_width7_depth9
  #(
    .init_file("./c_n.rom"),
    .read_f(1),
    .write_f(1),
    .output_file("./c_n_out.rom")
  )
  mem_2r_1w_width7_depth9
  (
    .clk(clk),
    .rd_addr0((rd)? rd_addr : { idx_in, ca_in }),
    .rd_addr1({ idx_in, cb_in }),
    .out0({ na_v_t, na_t }),
    .out1({ nb_v_t, nb_t }),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  fifo
  #(
    .FIFO_WIDTH(16),
    .FIFO_DEPTH_BITS(3)
  )
  fifo_a
  (
    .clk(clk),
    .rst(rst),
    .write_enable(fifoa_wr_en),
    .input_data(fifoa_data),
    .output_read_enable(fifoa_rd_en),
    .output_data(wa_t)
  );


  fifo
  #(
    .FIFO_WIDTH(16),
    .FIFO_DEPTH_BITS(3)
  )
  fifo_b
  (
    .clk(clk),
    .rst(rst),
    .write_enable(fifob_wr_en),
    .input_data(fifob_data),
    .output_read_enable(fifob_rd_en),
    .output_data(wb_t)
  );


  initial begin
    out_v = 0;
    out_data = 0;
    rdy = 0;
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    na_out = 0;
    na_v_out = 0;
    nb_out = 0;
    nb_v_out = 0;
    sw_out = 0;
    wa_out = 0;
    wb_out = 0;
    flag = 0;
    counter = 0;
    fifo_init = 0;
  end


endmodule



module mem_2r_1w_width7_depth9 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [9-1:0] rd_addr0,
  input [9-1:0] rd_addr1,
  output [7-1:0] out0,
  output [7-1:0] out1,
  input wr,
  input [9-1:0] wr_addr,
  input [7-1:0] wr_data
);

  (*rom_style = "block" *) reg [7-1:0] mem[0:2**9-1];
  /*
  reg [7-1:0] mem [0:2**9-1];
  */
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end

  //synthesis translate_on

  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end


endmodule



module fifo #
(
  parameter FIFO_WIDTH = 32,
  parameter FIFO_DEPTH_BITS = 8,
  parameter FIFO_ALMOSTFULL_THRESHOLD = 2 ** FIFO_DEPTH_BITS - 4,
  parameter FIFO_ALMOSTEMPTY_THRESHOLD = 4
)
(
  input clk,
  input rst,
  input write_enable,
  input [FIFO_WIDTH-1:0] input_data,
  input output_read_enable,
  output reg output_valid,
  output reg [FIFO_WIDTH-1:0] output_data,
  output reg empty,
  output reg almostempty,
  output reg full,
  output reg almostfull,
  output reg [FIFO_DEPTH_BITS+1-1:0] data_count
);

  reg [FIFO_DEPTH_BITS-1:0] read_pointer;
  reg [FIFO_DEPTH_BITS-1:0] write_pointer;
  (*rom_style = "block" *) reg [FIFO_WIDTH-1:0] mem[0:2**FIFO_DEPTH_BITS-1];
  /*
  reg [FIFO_WIDTH-1:0] mem [0:2**FIFO_DEPTH_BITS-1];
  */

  always @(posedge clk) begin
    if(rst) begin
      empty <= 1;
      almostempty <= 1;
      full <= 0;
      almostfull <= 0;
      read_pointer <= 0;
      write_pointer <= 0;
      data_count <= 0;
    end else begin
      case({ write_enable, output_read_enable })
        3: begin
          read_pointer <= read_pointer + 1;
          write_pointer <= write_pointer + 1;
        end
        2: begin
          if(~full) begin
            write_pointer <= write_pointer + 1;
            data_count <= data_count + 1;
            empty <= 0;
            if(data_count == FIFO_ALMOSTEMPTY_THRESHOLD - 1) begin
              almostempty <= 0;
            end 
            if(data_count == 2 ** FIFO_DEPTH_BITS - 1) begin
              full <= 1;
            end 
            if(data_count == FIFO_ALMOSTFULL_THRESHOLD - 1) begin
              almostfull <= 1;
            end 
          end 
        end
        1: begin
          if(~empty) begin
            read_pointer <= read_pointer + 1;
            data_count <= data_count - 1;
            full <= 0;
            if(data_count == FIFO_ALMOSTFULL_THRESHOLD) begin
              almostfull <= 0;
            end 
            if(data_count == 1) begin
              empty <= 1;
            end 
            if(data_count == FIFO_ALMOSTEMPTY_THRESHOLD) begin
              almostempty <= 1;
            end 
          end 
        end
      endcase
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      output_valid <= 0;
    end else begin
      output_valid <= 0;
      if(write_enable == 1) begin
        mem[write_pointer] <= input_data;
      end 
      if(output_read_enable == 1) begin
        output_data <= mem[read_pointer];
        output_valid <= 1;
      end 
    end
  end


endmodule



module st2_n_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [6-1:0] ca_in,
  input [6-1:0] cb_in,
  input [6-1:0] na_in,
  input na_v_in,
  input [6-1:0] nb_in,
  input nb_v_in,
  input sw_in,
  input [16-1:0] wa_in,
  input [16-1:0] wb_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [6-1:0] ca_out,
  output reg [6-1:0] cb_out,
  output reg [6-1:0] na_out,
  output reg na_v_out,
  output reg [6-1:0] nb_out,
  output reg nb_v_out,
  output reg [24-1:0] va_out,
  output reg [4-1:0] va_v_out,
  output reg [24-1:0] vb_out,
  output reg [4-1:0] vb_v_out,
  output reg sw_out,
  output reg [16-1:0] wa_out,
  output reg [16-1:0] wb_out
);

  wire [24-1:0] va_t;
  wire [4-1:0] va_v_t;
  wire [4-1:0] va_v_m;
  wire [24-1:0] vb_t;
  wire [4-1:0] vb_v_t;
  wire [4-1:0] vb_v_m;
  assign va_v_t = (na_v_in)? va_v_m : 4'b0;
  assign vb_v_t = (nb_v_in)? vb_v_m : 4'b0;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    na_out <= na_in;
    na_v_out <= na_v_in;
    nb_out <= nb_in;
    nb_v_out <= nb_v_in;
    sw_out <= sw_in;
    wa_out <= wa_in;
    wb_out <= wb_in;
    va_out <= va_t;
    va_v_out <= va_v_t;
    vb_out <= vb_t;
    vb_v_out <= vb_v_t;
  end


  mem_2r_1w_width7_depth6
  #(
    .init_file("./n0.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width7_depth6_0
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[0], va_t[5:0] }),
    .out1({ vb_v_m[0], vb_t[5:0] }),
    .wr(1'b0),
    .wr_addr(6'b0),
    .wr_data(7'b0)
  );


  mem_2r_1w_width7_depth6
  #(
    .init_file("./n1.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width7_depth6_1
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[1], va_t[11:6] }),
    .out1({ vb_v_m[1], vb_t[11:6] }),
    .wr(1'b0),
    .wr_addr(6'b0),
    .wr_data(7'b0)
  );


  mem_2r_1w_width7_depth6
  #(
    .init_file("./n2.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width7_depth6_2
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[2], va_t[17:12] }),
    .out1({ vb_v_m[2], vb_t[17:12] }),
    .wr(1'b0),
    .wr_addr(6'b0),
    .wr_data(7'b0)
  );


  mem_2r_1w_width7_depth6
  #(
    .init_file("./n3.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width7_depth6_3
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[3], va_t[23:18] }),
    .out1({ vb_v_m[3], vb_t[23:18] }),
    .wr(1'b0),
    .wr_addr(6'b0),
    .wr_data(7'b0)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    na_out = 0;
    na_v_out = 0;
    nb_out = 0;
    nb_v_out = 0;
    va_out = 0;
    va_v_out = 0;
    vb_out = 0;
    vb_v_out = 0;
    sw_out = 0;
    wa_out = 0;
    wb_out = 0;
  end


endmodule



module mem_2r_1w_width7_depth6 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [6-1:0] rd_addr0,
  input [6-1:0] rd_addr1,
  output [7-1:0] out0,
  output [7-1:0] out1,
  input wr,
  input [6-1:0] wr_addr,
  input [7-1:0] wr_data
);

  (*rom_style = "block" *) reg [7-1:0] mem[0:2**6-1];
  /*
  reg [7-1:0] mem [0:2**6-1];
  */
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end

  //synthesis translate_on

  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end


endmodule



module st3_n2c_6th_64cells
(
  input clk,
  input rst,
  input [3-1:0] idx_in,
  input v_in,
  input [6-1:0] ca_in,
  input [6-1:0] cb_in,
  input [6-1:0] na_in,
  input na_v_in,
  input [6-1:0] nb_in,
  input nb_v_in,
  input [24-1:0] va_in,
  input [4-1:0] va_v_in,
  input [24-1:0] vb_in,
  input [4-1:0] vb_v_in,
  input [16-1:0] st3_wb_in,
  input sw_in,
  input [16-1:0] wa_in,
  input [16-1:0] wb_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [6-1:0] ca_out,
  output reg [6-1:0] cb_out,
  output reg [24-1:0] cva_out,
  output reg [4-1:0] cva_v_out,
  output reg [24-1:0] cvb_out,
  output reg [4-1:0] cvb_v_out,
  output reg [16-1:0] wb_out
);

  reg flag;
  wire [24-1:0] cva_t;
  wire [24-1:0] cvb_t;
  wire [3-1:0] wa_idx;
  wire [6-1:0] wa_c;
  wire [6-1:0] wa_n;
  wire wa_n_v;
  wire [3-1:0] wb_idx;
  wire [6-1:0] wb_c;
  wire [6-1:0] wb_n;
  wire wb_n_v;
  wire m_wr;
  wire [9-1:0] m_wr_addr;
  wire [6-1:0] m_wr_data;
  assign wa_n = wa_in[5:0];
  assign wa_n_v = wa_in[6];
  assign wa_c = wa_in[12:7];
  assign wa_idx = wa_in[15:13];
  assign wb_n = st3_wb_in[5:0];
  assign wb_n_v = st3_wb_in[6];
  assign wb_c = st3_wb_in[12:7];
  assign wb_idx = st3_wb_in[15:13];
  assign m_wr = (flag)? &{ sw_in, wa_n_v } : &{ sw_in, wb_n_v };
  assign m_wr_addr = (flag)? { wa_idx, wa_n } : { wb_idx, wb_n };
  assign m_wr_data = (flag)? wa_c : wb_c;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    cva_out <= cva_t;
    cva_v_out <= va_v_in;
    cvb_out <= cvb_t;
    cvb_v_out <= vb_v_in;
    wb_out <= wb_in;
  end


  always @(posedge clk) begin
    if(rst) begin
      flag <= 1;
    end else begin
      if(sw_in) begin
        flag <= ~flag;
      end 
    end
  end


  mem_2r_1w_width6_depth9
  #(
    .init_file("./n_c.rom"),
    .read_f(1),
    .write_f(1),
    .output_file("./n_c_out.rom")
  )
  mem_2r_1w_width6_depth9_0
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[5:0] }),
    .rd_addr1({ idx_in, vb_in[5:0] }),
    .out0(cva_t[5:0]),
    .out1(cvb_t[5:0]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width6_depth9
  #(
    .init_file("./n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./n_c_out.rom")
  )
  mem_2r_1w_width6_depth9_1
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[11:6] }),
    .rd_addr1({ idx_in, vb_in[11:6] }),
    .out0(cva_t[11:6]),
    .out1(cvb_t[11:6]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width6_depth9
  #(
    .init_file("./n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./n_c_out.rom")
  )
  mem_2r_1w_width6_depth9_2
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[17:12] }),
    .rd_addr1({ idx_in, vb_in[17:12] }),
    .out0(cva_t[17:12]),
    .out1(cvb_t[17:12]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width6_depth9
  #(
    .init_file("./n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./n_c_out.rom")
  )
  mem_2r_1w_width6_depth9_3
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[23:18] }),
    .rd_addr1({ idx_in, vb_in[23:18] }),
    .out0(cva_t[23:18]),
    .out1(cvb_t[23:18]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    cva_out = 0;
    cva_v_out = 0;
    cvb_out = 0;
    cvb_v_out = 0;
    wb_out = 0;
    flag = 0;
  end


endmodule



module mem_2r_1w_width6_depth9 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [9-1:0] rd_addr0,
  input [9-1:0] rd_addr1,
  output [6-1:0] out0,
  output [6-1:0] out1,
  input wr,
  input [9-1:0] wr_addr,
  input [6-1:0] wr_data
);

  (*rom_style = "block" *) reg [6-1:0] mem[0:2**9-1];
  /*
  reg [6-1:0] mem [0:2**9-1];
  */
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end

  //synthesis translate_on

  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end


endmodule



module st4_d1_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [6-1:0] ca_in,
  input [6-1:0] cb_in,
  input [24-1:0] cva_in,
  input [4-1:0] cva_v_in,
  input [24-1:0] cvb_in,
  input [4-1:0] cvb_v_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [6-1:0] ca_out,
  output reg [6-1:0] cb_out,
  output reg [24-1:0] cva_out,
  output reg [4-1:0] cva_v_out,
  output reg [24-1:0] cvb_out,
  output reg [4-1:0] cvb_v_out,
  output reg [36-1:0] dvac_out,
  output reg [36-1:0] dvbc_out
);

  wire [6-1:0] cac;
  wire [6-1:0] cbc;
  wire [36-1:0] dvac_t;
  wire [36-1:0] dvbc_t;
  assign cac = ca_in;
  assign cbc = cb_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    cva_out <= cva_in;
    cva_v_out <= cva_v_in;
    cvb_out <= cvb_in;
    cvb_v_out <= cvb_v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
  end


  distance_rom_8_8
  distance_rom_8_8_dac_0
  (
    .opa0(cac),
    .opa1(cva_in[5:0]),
    .opav(cva_v_in[0]),
    .opb0(cac),
    .opb1(cva_in[11:6]),
    .opbv(cva_v_in[1]),
    .da(dvac_t[8:0]),
    .db(dvac_t[17:9])
  );


  distance_rom_8_8
  distance_rom_8_8_dac_1
  (
    .opa0(cac),
    .opa1(cva_in[17:12]),
    .opav(cva_v_in[2]),
    .opb0(cac),
    .opb1(cva_in[23:18]),
    .opbv(cva_v_in[3]),
    .da(dvac_t[26:18]),
    .db(dvac_t[35:27])
  );


  distance_rom_8_8
  distance_rom_8_8_dbc_0
  (
    .opa0(cbc),
    .opa1(cvb_in[5:0]),
    .opav(cvb_v_in[0]),
    .opb0(cbc),
    .opb1(cvb_in[11:6]),
    .opbv(cvb_v_in[1]),
    .da(dvbc_t[8:0]),
    .db(dvbc_t[17:9])
  );


  distance_rom_8_8
  distance_rom_8_8_dbc_1
  (
    .opa0(cbc),
    .opa1(cvb_in[17:12]),
    .opav(cvb_v_in[2]),
    .opb0(cbc),
    .opb1(cvb_in[23:18]),
    .opbv(cvb_v_in[3]),
    .da(dvbc_t[26:18]),
    .db(dvbc_t[35:27])
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    cva_out = 0;
    cva_v_out = 0;
    cvb_out = 0;
    cvb_v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
  end


endmodule



module distance_rom_8_8
(
  input [6-1:0] opa0,
  input [6-1:0] opa1,
  input opav,
  input [6-1:0] opb0,
  input [6-1:0] opb1,
  input opbv,
  output [9-1:0] da,
  output [9-1:0] db
);

  wire [9-1:0] mem [0:64**2-1];
  assign da = (opav)? mem[{ opa1, opa0 }] : 0;
  assign db = (opbv)? mem[{ opb1, opb0 }] : 0;
  assign mem[0] = 9'd0;
  assign mem[1] = 9'd1;
  assign mem[2] = 9'd2;
  assign mem[3] = 9'd3;
  assign mem[4] = 9'd4;
  assign mem[5] = 9'd5;
  assign mem[6] = 9'd6;
  assign mem[7] = 9'd7;
  assign mem[8] = 9'd1;
  assign mem[9] = 9'd2;
  assign mem[10] = 9'd3;
  assign mem[11] = 9'd4;
  assign mem[12] = 9'd5;
  assign mem[13] = 9'd6;
  assign mem[14] = 9'd7;
  assign mem[15] = 9'd8;
  assign mem[16] = 9'd2;
  assign mem[17] = 9'd3;
  assign mem[18] = 9'd4;
  assign mem[19] = 9'd5;
  assign mem[20] = 9'd6;
  assign mem[21] = 9'd7;
  assign mem[22] = 9'd8;
  assign mem[23] = 9'd9;
  assign mem[24] = 9'd3;
  assign mem[25] = 9'd4;
  assign mem[26] = 9'd5;
  assign mem[27] = 9'd6;
  assign mem[28] = 9'd7;
  assign mem[29] = 9'd8;
  assign mem[30] = 9'd9;
  assign mem[31] = 9'd10;
  assign mem[32] = 9'd4;
  assign mem[33] = 9'd5;
  assign mem[34] = 9'd6;
  assign mem[35] = 9'd7;
  assign mem[36] = 9'd8;
  assign mem[37] = 9'd9;
  assign mem[38] = 9'd10;
  assign mem[39] = 9'd11;
  assign mem[40] = 9'd5;
  assign mem[41] = 9'd6;
  assign mem[42] = 9'd7;
  assign mem[43] = 9'd8;
  assign mem[44] = 9'd9;
  assign mem[45] = 9'd10;
  assign mem[46] = 9'd11;
  assign mem[47] = 9'd12;
  assign mem[48] = 9'd6;
  assign mem[49] = 9'd7;
  assign mem[50] = 9'd8;
  assign mem[51] = 9'd9;
  assign mem[52] = 9'd10;
  assign mem[53] = 9'd11;
  assign mem[54] = 9'd12;
  assign mem[55] = 9'd13;
  assign mem[56] = 9'd7;
  assign mem[57] = 9'd8;
  assign mem[58] = 9'd9;
  assign mem[59] = 9'd10;
  assign mem[60] = 9'd11;
  assign mem[61] = 9'd12;
  assign mem[62] = 9'd13;
  assign mem[63] = 9'd14;
  assign mem[64] = 9'd1;
  assign mem[65] = 9'd0;
  assign mem[66] = 9'd1;
  assign mem[67] = 9'd2;
  assign mem[68] = 9'd3;
  assign mem[69] = 9'd4;
  assign mem[70] = 9'd5;
  assign mem[71] = 9'd6;
  assign mem[72] = 9'd2;
  assign mem[73] = 9'd1;
  assign mem[74] = 9'd2;
  assign mem[75] = 9'd3;
  assign mem[76] = 9'd4;
  assign mem[77] = 9'd5;
  assign mem[78] = 9'd6;
  assign mem[79] = 9'd7;
  assign mem[80] = 9'd3;
  assign mem[81] = 9'd2;
  assign mem[82] = 9'd3;
  assign mem[83] = 9'd4;
  assign mem[84] = 9'd5;
  assign mem[85] = 9'd6;
  assign mem[86] = 9'd7;
  assign mem[87] = 9'd8;
  assign mem[88] = 9'd4;
  assign mem[89] = 9'd3;
  assign mem[90] = 9'd4;
  assign mem[91] = 9'd5;
  assign mem[92] = 9'd6;
  assign mem[93] = 9'd7;
  assign mem[94] = 9'd8;
  assign mem[95] = 9'd9;
  assign mem[96] = 9'd5;
  assign mem[97] = 9'd4;
  assign mem[98] = 9'd5;
  assign mem[99] = 9'd6;
  assign mem[100] = 9'd7;
  assign mem[101] = 9'd8;
  assign mem[102] = 9'd9;
  assign mem[103] = 9'd10;
  assign mem[104] = 9'd6;
  assign mem[105] = 9'd5;
  assign mem[106] = 9'd6;
  assign mem[107] = 9'd7;
  assign mem[108] = 9'd8;
  assign mem[109] = 9'd9;
  assign mem[110] = 9'd10;
  assign mem[111] = 9'd11;
  assign mem[112] = 9'd7;
  assign mem[113] = 9'd6;
  assign mem[114] = 9'd7;
  assign mem[115] = 9'd8;
  assign mem[116] = 9'd9;
  assign mem[117] = 9'd10;
  assign mem[118] = 9'd11;
  assign mem[119] = 9'd12;
  assign mem[120] = 9'd8;
  assign mem[121] = 9'd7;
  assign mem[122] = 9'd8;
  assign mem[123] = 9'd9;
  assign mem[124] = 9'd10;
  assign mem[125] = 9'd11;
  assign mem[126] = 9'd12;
  assign mem[127] = 9'd13;
  assign mem[128] = 9'd2;
  assign mem[129] = 9'd1;
  assign mem[130] = 9'd0;
  assign mem[131] = 9'd1;
  assign mem[132] = 9'd2;
  assign mem[133] = 9'd3;
  assign mem[134] = 9'd4;
  assign mem[135] = 9'd5;
  assign mem[136] = 9'd3;
  assign mem[137] = 9'd2;
  assign mem[138] = 9'd1;
  assign mem[139] = 9'd2;
  assign mem[140] = 9'd3;
  assign mem[141] = 9'd4;
  assign mem[142] = 9'd5;
  assign mem[143] = 9'd6;
  assign mem[144] = 9'd4;
  assign mem[145] = 9'd3;
  assign mem[146] = 9'd2;
  assign mem[147] = 9'd3;
  assign mem[148] = 9'd4;
  assign mem[149] = 9'd5;
  assign mem[150] = 9'd6;
  assign mem[151] = 9'd7;
  assign mem[152] = 9'd5;
  assign mem[153] = 9'd4;
  assign mem[154] = 9'd3;
  assign mem[155] = 9'd4;
  assign mem[156] = 9'd5;
  assign mem[157] = 9'd6;
  assign mem[158] = 9'd7;
  assign mem[159] = 9'd8;
  assign mem[160] = 9'd6;
  assign mem[161] = 9'd5;
  assign mem[162] = 9'd4;
  assign mem[163] = 9'd5;
  assign mem[164] = 9'd6;
  assign mem[165] = 9'd7;
  assign mem[166] = 9'd8;
  assign mem[167] = 9'd9;
  assign mem[168] = 9'd7;
  assign mem[169] = 9'd6;
  assign mem[170] = 9'd5;
  assign mem[171] = 9'd6;
  assign mem[172] = 9'd7;
  assign mem[173] = 9'd8;
  assign mem[174] = 9'd9;
  assign mem[175] = 9'd10;
  assign mem[176] = 9'd8;
  assign mem[177] = 9'd7;
  assign mem[178] = 9'd6;
  assign mem[179] = 9'd7;
  assign mem[180] = 9'd8;
  assign mem[181] = 9'd9;
  assign mem[182] = 9'd10;
  assign mem[183] = 9'd11;
  assign mem[184] = 9'd9;
  assign mem[185] = 9'd8;
  assign mem[186] = 9'd7;
  assign mem[187] = 9'd8;
  assign mem[188] = 9'd9;
  assign mem[189] = 9'd10;
  assign mem[190] = 9'd11;
  assign mem[191] = 9'd12;
  assign mem[192] = 9'd3;
  assign mem[193] = 9'd2;
  assign mem[194] = 9'd1;
  assign mem[195] = 9'd0;
  assign mem[196] = 9'd1;
  assign mem[197] = 9'd2;
  assign mem[198] = 9'd3;
  assign mem[199] = 9'd4;
  assign mem[200] = 9'd4;
  assign mem[201] = 9'd3;
  assign mem[202] = 9'd2;
  assign mem[203] = 9'd1;
  assign mem[204] = 9'd2;
  assign mem[205] = 9'd3;
  assign mem[206] = 9'd4;
  assign mem[207] = 9'd5;
  assign mem[208] = 9'd5;
  assign mem[209] = 9'd4;
  assign mem[210] = 9'd3;
  assign mem[211] = 9'd2;
  assign mem[212] = 9'd3;
  assign mem[213] = 9'd4;
  assign mem[214] = 9'd5;
  assign mem[215] = 9'd6;
  assign mem[216] = 9'd6;
  assign mem[217] = 9'd5;
  assign mem[218] = 9'd4;
  assign mem[219] = 9'd3;
  assign mem[220] = 9'd4;
  assign mem[221] = 9'd5;
  assign mem[222] = 9'd6;
  assign mem[223] = 9'd7;
  assign mem[224] = 9'd7;
  assign mem[225] = 9'd6;
  assign mem[226] = 9'd5;
  assign mem[227] = 9'd4;
  assign mem[228] = 9'd5;
  assign mem[229] = 9'd6;
  assign mem[230] = 9'd7;
  assign mem[231] = 9'd8;
  assign mem[232] = 9'd8;
  assign mem[233] = 9'd7;
  assign mem[234] = 9'd6;
  assign mem[235] = 9'd5;
  assign mem[236] = 9'd6;
  assign mem[237] = 9'd7;
  assign mem[238] = 9'd8;
  assign mem[239] = 9'd9;
  assign mem[240] = 9'd9;
  assign mem[241] = 9'd8;
  assign mem[242] = 9'd7;
  assign mem[243] = 9'd6;
  assign mem[244] = 9'd7;
  assign mem[245] = 9'd8;
  assign mem[246] = 9'd9;
  assign mem[247] = 9'd10;
  assign mem[248] = 9'd10;
  assign mem[249] = 9'd9;
  assign mem[250] = 9'd8;
  assign mem[251] = 9'd7;
  assign mem[252] = 9'd8;
  assign mem[253] = 9'd9;
  assign mem[254] = 9'd10;
  assign mem[255] = 9'd11;
  assign mem[256] = 9'd4;
  assign mem[257] = 9'd3;
  assign mem[258] = 9'd2;
  assign mem[259] = 9'd1;
  assign mem[260] = 9'd0;
  assign mem[261] = 9'd1;
  assign mem[262] = 9'd2;
  assign mem[263] = 9'd3;
  assign mem[264] = 9'd5;
  assign mem[265] = 9'd4;
  assign mem[266] = 9'd3;
  assign mem[267] = 9'd2;
  assign mem[268] = 9'd1;
  assign mem[269] = 9'd2;
  assign mem[270] = 9'd3;
  assign mem[271] = 9'd4;
  assign mem[272] = 9'd6;
  assign mem[273] = 9'd5;
  assign mem[274] = 9'd4;
  assign mem[275] = 9'd3;
  assign mem[276] = 9'd2;
  assign mem[277] = 9'd3;
  assign mem[278] = 9'd4;
  assign mem[279] = 9'd5;
  assign mem[280] = 9'd7;
  assign mem[281] = 9'd6;
  assign mem[282] = 9'd5;
  assign mem[283] = 9'd4;
  assign mem[284] = 9'd3;
  assign mem[285] = 9'd4;
  assign mem[286] = 9'd5;
  assign mem[287] = 9'd6;
  assign mem[288] = 9'd8;
  assign mem[289] = 9'd7;
  assign mem[290] = 9'd6;
  assign mem[291] = 9'd5;
  assign mem[292] = 9'd4;
  assign mem[293] = 9'd5;
  assign mem[294] = 9'd6;
  assign mem[295] = 9'd7;
  assign mem[296] = 9'd9;
  assign mem[297] = 9'd8;
  assign mem[298] = 9'd7;
  assign mem[299] = 9'd6;
  assign mem[300] = 9'd5;
  assign mem[301] = 9'd6;
  assign mem[302] = 9'd7;
  assign mem[303] = 9'd8;
  assign mem[304] = 9'd10;
  assign mem[305] = 9'd9;
  assign mem[306] = 9'd8;
  assign mem[307] = 9'd7;
  assign mem[308] = 9'd6;
  assign mem[309] = 9'd7;
  assign mem[310] = 9'd8;
  assign mem[311] = 9'd9;
  assign mem[312] = 9'd11;
  assign mem[313] = 9'd10;
  assign mem[314] = 9'd9;
  assign mem[315] = 9'd8;
  assign mem[316] = 9'd7;
  assign mem[317] = 9'd8;
  assign mem[318] = 9'd9;
  assign mem[319] = 9'd10;
  assign mem[320] = 9'd5;
  assign mem[321] = 9'd4;
  assign mem[322] = 9'd3;
  assign mem[323] = 9'd2;
  assign mem[324] = 9'd1;
  assign mem[325] = 9'd0;
  assign mem[326] = 9'd1;
  assign mem[327] = 9'd2;
  assign mem[328] = 9'd6;
  assign mem[329] = 9'd5;
  assign mem[330] = 9'd4;
  assign mem[331] = 9'd3;
  assign mem[332] = 9'd2;
  assign mem[333] = 9'd1;
  assign mem[334] = 9'd2;
  assign mem[335] = 9'd3;
  assign mem[336] = 9'd7;
  assign mem[337] = 9'd6;
  assign mem[338] = 9'd5;
  assign mem[339] = 9'd4;
  assign mem[340] = 9'd3;
  assign mem[341] = 9'd2;
  assign mem[342] = 9'd3;
  assign mem[343] = 9'd4;
  assign mem[344] = 9'd8;
  assign mem[345] = 9'd7;
  assign mem[346] = 9'd6;
  assign mem[347] = 9'd5;
  assign mem[348] = 9'd4;
  assign mem[349] = 9'd3;
  assign mem[350] = 9'd4;
  assign mem[351] = 9'd5;
  assign mem[352] = 9'd9;
  assign mem[353] = 9'd8;
  assign mem[354] = 9'd7;
  assign mem[355] = 9'd6;
  assign mem[356] = 9'd5;
  assign mem[357] = 9'd4;
  assign mem[358] = 9'd5;
  assign mem[359] = 9'd6;
  assign mem[360] = 9'd10;
  assign mem[361] = 9'd9;
  assign mem[362] = 9'd8;
  assign mem[363] = 9'd7;
  assign mem[364] = 9'd6;
  assign mem[365] = 9'd5;
  assign mem[366] = 9'd6;
  assign mem[367] = 9'd7;
  assign mem[368] = 9'd11;
  assign mem[369] = 9'd10;
  assign mem[370] = 9'd9;
  assign mem[371] = 9'd8;
  assign mem[372] = 9'd7;
  assign mem[373] = 9'd6;
  assign mem[374] = 9'd7;
  assign mem[375] = 9'd8;
  assign mem[376] = 9'd12;
  assign mem[377] = 9'd11;
  assign mem[378] = 9'd10;
  assign mem[379] = 9'd9;
  assign mem[380] = 9'd8;
  assign mem[381] = 9'd7;
  assign mem[382] = 9'd8;
  assign mem[383] = 9'd9;
  assign mem[384] = 9'd6;
  assign mem[385] = 9'd5;
  assign mem[386] = 9'd4;
  assign mem[387] = 9'd3;
  assign mem[388] = 9'd2;
  assign mem[389] = 9'd1;
  assign mem[390] = 9'd0;
  assign mem[391] = 9'd1;
  assign mem[392] = 9'd7;
  assign mem[393] = 9'd6;
  assign mem[394] = 9'd5;
  assign mem[395] = 9'd4;
  assign mem[396] = 9'd3;
  assign mem[397] = 9'd2;
  assign mem[398] = 9'd1;
  assign mem[399] = 9'd2;
  assign mem[400] = 9'd8;
  assign mem[401] = 9'd7;
  assign mem[402] = 9'd6;
  assign mem[403] = 9'd5;
  assign mem[404] = 9'd4;
  assign mem[405] = 9'd3;
  assign mem[406] = 9'd2;
  assign mem[407] = 9'd3;
  assign mem[408] = 9'd9;
  assign mem[409] = 9'd8;
  assign mem[410] = 9'd7;
  assign mem[411] = 9'd6;
  assign mem[412] = 9'd5;
  assign mem[413] = 9'd4;
  assign mem[414] = 9'd3;
  assign mem[415] = 9'd4;
  assign mem[416] = 9'd10;
  assign mem[417] = 9'd9;
  assign mem[418] = 9'd8;
  assign mem[419] = 9'd7;
  assign mem[420] = 9'd6;
  assign mem[421] = 9'd5;
  assign mem[422] = 9'd4;
  assign mem[423] = 9'd5;
  assign mem[424] = 9'd11;
  assign mem[425] = 9'd10;
  assign mem[426] = 9'd9;
  assign mem[427] = 9'd8;
  assign mem[428] = 9'd7;
  assign mem[429] = 9'd6;
  assign mem[430] = 9'd5;
  assign mem[431] = 9'd6;
  assign mem[432] = 9'd12;
  assign mem[433] = 9'd11;
  assign mem[434] = 9'd10;
  assign mem[435] = 9'd9;
  assign mem[436] = 9'd8;
  assign mem[437] = 9'd7;
  assign mem[438] = 9'd6;
  assign mem[439] = 9'd7;
  assign mem[440] = 9'd13;
  assign mem[441] = 9'd12;
  assign mem[442] = 9'd11;
  assign mem[443] = 9'd10;
  assign mem[444] = 9'd9;
  assign mem[445] = 9'd8;
  assign mem[446] = 9'd7;
  assign mem[447] = 9'd8;
  assign mem[448] = 9'd7;
  assign mem[449] = 9'd6;
  assign mem[450] = 9'd5;
  assign mem[451] = 9'd4;
  assign mem[452] = 9'd3;
  assign mem[453] = 9'd2;
  assign mem[454] = 9'd1;
  assign mem[455] = 9'd0;
  assign mem[456] = 9'd8;
  assign mem[457] = 9'd7;
  assign mem[458] = 9'd6;
  assign mem[459] = 9'd5;
  assign mem[460] = 9'd4;
  assign mem[461] = 9'd3;
  assign mem[462] = 9'd2;
  assign mem[463] = 9'd1;
  assign mem[464] = 9'd9;
  assign mem[465] = 9'd8;
  assign mem[466] = 9'd7;
  assign mem[467] = 9'd6;
  assign mem[468] = 9'd5;
  assign mem[469] = 9'd4;
  assign mem[470] = 9'd3;
  assign mem[471] = 9'd2;
  assign mem[472] = 9'd10;
  assign mem[473] = 9'd9;
  assign mem[474] = 9'd8;
  assign mem[475] = 9'd7;
  assign mem[476] = 9'd6;
  assign mem[477] = 9'd5;
  assign mem[478] = 9'd4;
  assign mem[479] = 9'd3;
  assign mem[480] = 9'd11;
  assign mem[481] = 9'd10;
  assign mem[482] = 9'd9;
  assign mem[483] = 9'd8;
  assign mem[484] = 9'd7;
  assign mem[485] = 9'd6;
  assign mem[486] = 9'd5;
  assign mem[487] = 9'd4;
  assign mem[488] = 9'd12;
  assign mem[489] = 9'd11;
  assign mem[490] = 9'd10;
  assign mem[491] = 9'd9;
  assign mem[492] = 9'd8;
  assign mem[493] = 9'd7;
  assign mem[494] = 9'd6;
  assign mem[495] = 9'd5;
  assign mem[496] = 9'd13;
  assign mem[497] = 9'd12;
  assign mem[498] = 9'd11;
  assign mem[499] = 9'd10;
  assign mem[500] = 9'd9;
  assign mem[501] = 9'd8;
  assign mem[502] = 9'd7;
  assign mem[503] = 9'd6;
  assign mem[504] = 9'd14;
  assign mem[505] = 9'd13;
  assign mem[506] = 9'd12;
  assign mem[507] = 9'd11;
  assign mem[508] = 9'd10;
  assign mem[509] = 9'd9;
  assign mem[510] = 9'd8;
  assign mem[511] = 9'd7;
  assign mem[512] = 9'd1;
  assign mem[513] = 9'd2;
  assign mem[514] = 9'd3;
  assign mem[515] = 9'd4;
  assign mem[516] = 9'd5;
  assign mem[517] = 9'd6;
  assign mem[518] = 9'd7;
  assign mem[519] = 9'd8;
  assign mem[520] = 9'd0;
  assign mem[521] = 9'd1;
  assign mem[522] = 9'd2;
  assign mem[523] = 9'd3;
  assign mem[524] = 9'd4;
  assign mem[525] = 9'd5;
  assign mem[526] = 9'd6;
  assign mem[527] = 9'd7;
  assign mem[528] = 9'd1;
  assign mem[529] = 9'd2;
  assign mem[530] = 9'd3;
  assign mem[531] = 9'd4;
  assign mem[532] = 9'd5;
  assign mem[533] = 9'd6;
  assign mem[534] = 9'd7;
  assign mem[535] = 9'd8;
  assign mem[536] = 9'd2;
  assign mem[537] = 9'd3;
  assign mem[538] = 9'd4;
  assign mem[539] = 9'd5;
  assign mem[540] = 9'd6;
  assign mem[541] = 9'd7;
  assign mem[542] = 9'd8;
  assign mem[543] = 9'd9;
  assign mem[544] = 9'd3;
  assign mem[545] = 9'd4;
  assign mem[546] = 9'd5;
  assign mem[547] = 9'd6;
  assign mem[548] = 9'd7;
  assign mem[549] = 9'd8;
  assign mem[550] = 9'd9;
  assign mem[551] = 9'd10;
  assign mem[552] = 9'd4;
  assign mem[553] = 9'd5;
  assign mem[554] = 9'd6;
  assign mem[555] = 9'd7;
  assign mem[556] = 9'd8;
  assign mem[557] = 9'd9;
  assign mem[558] = 9'd10;
  assign mem[559] = 9'd11;
  assign mem[560] = 9'd5;
  assign mem[561] = 9'd6;
  assign mem[562] = 9'd7;
  assign mem[563] = 9'd8;
  assign mem[564] = 9'd9;
  assign mem[565] = 9'd10;
  assign mem[566] = 9'd11;
  assign mem[567] = 9'd12;
  assign mem[568] = 9'd6;
  assign mem[569] = 9'd7;
  assign mem[570] = 9'd8;
  assign mem[571] = 9'd9;
  assign mem[572] = 9'd10;
  assign mem[573] = 9'd11;
  assign mem[574] = 9'd12;
  assign mem[575] = 9'd13;
  assign mem[576] = 9'd2;
  assign mem[577] = 9'd1;
  assign mem[578] = 9'd2;
  assign mem[579] = 9'd3;
  assign mem[580] = 9'd4;
  assign mem[581] = 9'd5;
  assign mem[582] = 9'd6;
  assign mem[583] = 9'd7;
  assign mem[584] = 9'd1;
  assign mem[585] = 9'd0;
  assign mem[586] = 9'd1;
  assign mem[587] = 9'd2;
  assign mem[588] = 9'd3;
  assign mem[589] = 9'd4;
  assign mem[590] = 9'd5;
  assign mem[591] = 9'd6;
  assign mem[592] = 9'd2;
  assign mem[593] = 9'd1;
  assign mem[594] = 9'd2;
  assign mem[595] = 9'd3;
  assign mem[596] = 9'd4;
  assign mem[597] = 9'd5;
  assign mem[598] = 9'd6;
  assign mem[599] = 9'd7;
  assign mem[600] = 9'd3;
  assign mem[601] = 9'd2;
  assign mem[602] = 9'd3;
  assign mem[603] = 9'd4;
  assign mem[604] = 9'd5;
  assign mem[605] = 9'd6;
  assign mem[606] = 9'd7;
  assign mem[607] = 9'd8;
  assign mem[608] = 9'd4;
  assign mem[609] = 9'd3;
  assign mem[610] = 9'd4;
  assign mem[611] = 9'd5;
  assign mem[612] = 9'd6;
  assign mem[613] = 9'd7;
  assign mem[614] = 9'd8;
  assign mem[615] = 9'd9;
  assign mem[616] = 9'd5;
  assign mem[617] = 9'd4;
  assign mem[618] = 9'd5;
  assign mem[619] = 9'd6;
  assign mem[620] = 9'd7;
  assign mem[621] = 9'd8;
  assign mem[622] = 9'd9;
  assign mem[623] = 9'd10;
  assign mem[624] = 9'd6;
  assign mem[625] = 9'd5;
  assign mem[626] = 9'd6;
  assign mem[627] = 9'd7;
  assign mem[628] = 9'd8;
  assign mem[629] = 9'd9;
  assign mem[630] = 9'd10;
  assign mem[631] = 9'd11;
  assign mem[632] = 9'd7;
  assign mem[633] = 9'd6;
  assign mem[634] = 9'd7;
  assign mem[635] = 9'd8;
  assign mem[636] = 9'd9;
  assign mem[637] = 9'd10;
  assign mem[638] = 9'd11;
  assign mem[639] = 9'd12;
  assign mem[640] = 9'd3;
  assign mem[641] = 9'd2;
  assign mem[642] = 9'd1;
  assign mem[643] = 9'd2;
  assign mem[644] = 9'd3;
  assign mem[645] = 9'd4;
  assign mem[646] = 9'd5;
  assign mem[647] = 9'd6;
  assign mem[648] = 9'd2;
  assign mem[649] = 9'd1;
  assign mem[650] = 9'd0;
  assign mem[651] = 9'd1;
  assign mem[652] = 9'd2;
  assign mem[653] = 9'd3;
  assign mem[654] = 9'd4;
  assign mem[655] = 9'd5;
  assign mem[656] = 9'd3;
  assign mem[657] = 9'd2;
  assign mem[658] = 9'd1;
  assign mem[659] = 9'd2;
  assign mem[660] = 9'd3;
  assign mem[661] = 9'd4;
  assign mem[662] = 9'd5;
  assign mem[663] = 9'd6;
  assign mem[664] = 9'd4;
  assign mem[665] = 9'd3;
  assign mem[666] = 9'd2;
  assign mem[667] = 9'd3;
  assign mem[668] = 9'd4;
  assign mem[669] = 9'd5;
  assign mem[670] = 9'd6;
  assign mem[671] = 9'd7;
  assign mem[672] = 9'd5;
  assign mem[673] = 9'd4;
  assign mem[674] = 9'd3;
  assign mem[675] = 9'd4;
  assign mem[676] = 9'd5;
  assign mem[677] = 9'd6;
  assign mem[678] = 9'd7;
  assign mem[679] = 9'd8;
  assign mem[680] = 9'd6;
  assign mem[681] = 9'd5;
  assign mem[682] = 9'd4;
  assign mem[683] = 9'd5;
  assign mem[684] = 9'd6;
  assign mem[685] = 9'd7;
  assign mem[686] = 9'd8;
  assign mem[687] = 9'd9;
  assign mem[688] = 9'd7;
  assign mem[689] = 9'd6;
  assign mem[690] = 9'd5;
  assign mem[691] = 9'd6;
  assign mem[692] = 9'd7;
  assign mem[693] = 9'd8;
  assign mem[694] = 9'd9;
  assign mem[695] = 9'd10;
  assign mem[696] = 9'd8;
  assign mem[697] = 9'd7;
  assign mem[698] = 9'd6;
  assign mem[699] = 9'd7;
  assign mem[700] = 9'd8;
  assign mem[701] = 9'd9;
  assign mem[702] = 9'd10;
  assign mem[703] = 9'd11;
  assign mem[704] = 9'd4;
  assign mem[705] = 9'd3;
  assign mem[706] = 9'd2;
  assign mem[707] = 9'd1;
  assign mem[708] = 9'd2;
  assign mem[709] = 9'd3;
  assign mem[710] = 9'd4;
  assign mem[711] = 9'd5;
  assign mem[712] = 9'd3;
  assign mem[713] = 9'd2;
  assign mem[714] = 9'd1;
  assign mem[715] = 9'd0;
  assign mem[716] = 9'd1;
  assign mem[717] = 9'd2;
  assign mem[718] = 9'd3;
  assign mem[719] = 9'd4;
  assign mem[720] = 9'd4;
  assign mem[721] = 9'd3;
  assign mem[722] = 9'd2;
  assign mem[723] = 9'd1;
  assign mem[724] = 9'd2;
  assign mem[725] = 9'd3;
  assign mem[726] = 9'd4;
  assign mem[727] = 9'd5;
  assign mem[728] = 9'd5;
  assign mem[729] = 9'd4;
  assign mem[730] = 9'd3;
  assign mem[731] = 9'd2;
  assign mem[732] = 9'd3;
  assign mem[733] = 9'd4;
  assign mem[734] = 9'd5;
  assign mem[735] = 9'd6;
  assign mem[736] = 9'd6;
  assign mem[737] = 9'd5;
  assign mem[738] = 9'd4;
  assign mem[739] = 9'd3;
  assign mem[740] = 9'd4;
  assign mem[741] = 9'd5;
  assign mem[742] = 9'd6;
  assign mem[743] = 9'd7;
  assign mem[744] = 9'd7;
  assign mem[745] = 9'd6;
  assign mem[746] = 9'd5;
  assign mem[747] = 9'd4;
  assign mem[748] = 9'd5;
  assign mem[749] = 9'd6;
  assign mem[750] = 9'd7;
  assign mem[751] = 9'd8;
  assign mem[752] = 9'd8;
  assign mem[753] = 9'd7;
  assign mem[754] = 9'd6;
  assign mem[755] = 9'd5;
  assign mem[756] = 9'd6;
  assign mem[757] = 9'd7;
  assign mem[758] = 9'd8;
  assign mem[759] = 9'd9;
  assign mem[760] = 9'd9;
  assign mem[761] = 9'd8;
  assign mem[762] = 9'd7;
  assign mem[763] = 9'd6;
  assign mem[764] = 9'd7;
  assign mem[765] = 9'd8;
  assign mem[766] = 9'd9;
  assign mem[767] = 9'd10;
  assign mem[768] = 9'd5;
  assign mem[769] = 9'd4;
  assign mem[770] = 9'd3;
  assign mem[771] = 9'd2;
  assign mem[772] = 9'd1;
  assign mem[773] = 9'd2;
  assign mem[774] = 9'd3;
  assign mem[775] = 9'd4;
  assign mem[776] = 9'd4;
  assign mem[777] = 9'd3;
  assign mem[778] = 9'd2;
  assign mem[779] = 9'd1;
  assign mem[780] = 9'd0;
  assign mem[781] = 9'd1;
  assign mem[782] = 9'd2;
  assign mem[783] = 9'd3;
  assign mem[784] = 9'd5;
  assign mem[785] = 9'd4;
  assign mem[786] = 9'd3;
  assign mem[787] = 9'd2;
  assign mem[788] = 9'd1;
  assign mem[789] = 9'd2;
  assign mem[790] = 9'd3;
  assign mem[791] = 9'd4;
  assign mem[792] = 9'd6;
  assign mem[793] = 9'd5;
  assign mem[794] = 9'd4;
  assign mem[795] = 9'd3;
  assign mem[796] = 9'd2;
  assign mem[797] = 9'd3;
  assign mem[798] = 9'd4;
  assign mem[799] = 9'd5;
  assign mem[800] = 9'd7;
  assign mem[801] = 9'd6;
  assign mem[802] = 9'd5;
  assign mem[803] = 9'd4;
  assign mem[804] = 9'd3;
  assign mem[805] = 9'd4;
  assign mem[806] = 9'd5;
  assign mem[807] = 9'd6;
  assign mem[808] = 9'd8;
  assign mem[809] = 9'd7;
  assign mem[810] = 9'd6;
  assign mem[811] = 9'd5;
  assign mem[812] = 9'd4;
  assign mem[813] = 9'd5;
  assign mem[814] = 9'd6;
  assign mem[815] = 9'd7;
  assign mem[816] = 9'd9;
  assign mem[817] = 9'd8;
  assign mem[818] = 9'd7;
  assign mem[819] = 9'd6;
  assign mem[820] = 9'd5;
  assign mem[821] = 9'd6;
  assign mem[822] = 9'd7;
  assign mem[823] = 9'd8;
  assign mem[824] = 9'd10;
  assign mem[825] = 9'd9;
  assign mem[826] = 9'd8;
  assign mem[827] = 9'd7;
  assign mem[828] = 9'd6;
  assign mem[829] = 9'd7;
  assign mem[830] = 9'd8;
  assign mem[831] = 9'd9;
  assign mem[832] = 9'd6;
  assign mem[833] = 9'd5;
  assign mem[834] = 9'd4;
  assign mem[835] = 9'd3;
  assign mem[836] = 9'd2;
  assign mem[837] = 9'd1;
  assign mem[838] = 9'd2;
  assign mem[839] = 9'd3;
  assign mem[840] = 9'd5;
  assign mem[841] = 9'd4;
  assign mem[842] = 9'd3;
  assign mem[843] = 9'd2;
  assign mem[844] = 9'd1;
  assign mem[845] = 9'd0;
  assign mem[846] = 9'd1;
  assign mem[847] = 9'd2;
  assign mem[848] = 9'd6;
  assign mem[849] = 9'd5;
  assign mem[850] = 9'd4;
  assign mem[851] = 9'd3;
  assign mem[852] = 9'd2;
  assign mem[853] = 9'd1;
  assign mem[854] = 9'd2;
  assign mem[855] = 9'd3;
  assign mem[856] = 9'd7;
  assign mem[857] = 9'd6;
  assign mem[858] = 9'd5;
  assign mem[859] = 9'd4;
  assign mem[860] = 9'd3;
  assign mem[861] = 9'd2;
  assign mem[862] = 9'd3;
  assign mem[863] = 9'd4;
  assign mem[864] = 9'd8;
  assign mem[865] = 9'd7;
  assign mem[866] = 9'd6;
  assign mem[867] = 9'd5;
  assign mem[868] = 9'd4;
  assign mem[869] = 9'd3;
  assign mem[870] = 9'd4;
  assign mem[871] = 9'd5;
  assign mem[872] = 9'd9;
  assign mem[873] = 9'd8;
  assign mem[874] = 9'd7;
  assign mem[875] = 9'd6;
  assign mem[876] = 9'd5;
  assign mem[877] = 9'd4;
  assign mem[878] = 9'd5;
  assign mem[879] = 9'd6;
  assign mem[880] = 9'd10;
  assign mem[881] = 9'd9;
  assign mem[882] = 9'd8;
  assign mem[883] = 9'd7;
  assign mem[884] = 9'd6;
  assign mem[885] = 9'd5;
  assign mem[886] = 9'd6;
  assign mem[887] = 9'd7;
  assign mem[888] = 9'd11;
  assign mem[889] = 9'd10;
  assign mem[890] = 9'd9;
  assign mem[891] = 9'd8;
  assign mem[892] = 9'd7;
  assign mem[893] = 9'd6;
  assign mem[894] = 9'd7;
  assign mem[895] = 9'd8;
  assign mem[896] = 9'd7;
  assign mem[897] = 9'd6;
  assign mem[898] = 9'd5;
  assign mem[899] = 9'd4;
  assign mem[900] = 9'd3;
  assign mem[901] = 9'd2;
  assign mem[902] = 9'd1;
  assign mem[903] = 9'd2;
  assign mem[904] = 9'd6;
  assign mem[905] = 9'd5;
  assign mem[906] = 9'd4;
  assign mem[907] = 9'd3;
  assign mem[908] = 9'd2;
  assign mem[909] = 9'd1;
  assign mem[910] = 9'd0;
  assign mem[911] = 9'd1;
  assign mem[912] = 9'd7;
  assign mem[913] = 9'd6;
  assign mem[914] = 9'd5;
  assign mem[915] = 9'd4;
  assign mem[916] = 9'd3;
  assign mem[917] = 9'd2;
  assign mem[918] = 9'd1;
  assign mem[919] = 9'd2;
  assign mem[920] = 9'd8;
  assign mem[921] = 9'd7;
  assign mem[922] = 9'd6;
  assign mem[923] = 9'd5;
  assign mem[924] = 9'd4;
  assign mem[925] = 9'd3;
  assign mem[926] = 9'd2;
  assign mem[927] = 9'd3;
  assign mem[928] = 9'd9;
  assign mem[929] = 9'd8;
  assign mem[930] = 9'd7;
  assign mem[931] = 9'd6;
  assign mem[932] = 9'd5;
  assign mem[933] = 9'd4;
  assign mem[934] = 9'd3;
  assign mem[935] = 9'd4;
  assign mem[936] = 9'd10;
  assign mem[937] = 9'd9;
  assign mem[938] = 9'd8;
  assign mem[939] = 9'd7;
  assign mem[940] = 9'd6;
  assign mem[941] = 9'd5;
  assign mem[942] = 9'd4;
  assign mem[943] = 9'd5;
  assign mem[944] = 9'd11;
  assign mem[945] = 9'd10;
  assign mem[946] = 9'd9;
  assign mem[947] = 9'd8;
  assign mem[948] = 9'd7;
  assign mem[949] = 9'd6;
  assign mem[950] = 9'd5;
  assign mem[951] = 9'd6;
  assign mem[952] = 9'd12;
  assign mem[953] = 9'd11;
  assign mem[954] = 9'd10;
  assign mem[955] = 9'd9;
  assign mem[956] = 9'd8;
  assign mem[957] = 9'd7;
  assign mem[958] = 9'd6;
  assign mem[959] = 9'd7;
  assign mem[960] = 9'd8;
  assign mem[961] = 9'd7;
  assign mem[962] = 9'd6;
  assign mem[963] = 9'd5;
  assign mem[964] = 9'd4;
  assign mem[965] = 9'd3;
  assign mem[966] = 9'd2;
  assign mem[967] = 9'd1;
  assign mem[968] = 9'd7;
  assign mem[969] = 9'd6;
  assign mem[970] = 9'd5;
  assign mem[971] = 9'd4;
  assign mem[972] = 9'd3;
  assign mem[973] = 9'd2;
  assign mem[974] = 9'd1;
  assign mem[975] = 9'd0;
  assign mem[976] = 9'd8;
  assign mem[977] = 9'd7;
  assign mem[978] = 9'd6;
  assign mem[979] = 9'd5;
  assign mem[980] = 9'd4;
  assign mem[981] = 9'd3;
  assign mem[982] = 9'd2;
  assign mem[983] = 9'd1;
  assign mem[984] = 9'd9;
  assign mem[985] = 9'd8;
  assign mem[986] = 9'd7;
  assign mem[987] = 9'd6;
  assign mem[988] = 9'd5;
  assign mem[989] = 9'd4;
  assign mem[990] = 9'd3;
  assign mem[991] = 9'd2;
  assign mem[992] = 9'd10;
  assign mem[993] = 9'd9;
  assign mem[994] = 9'd8;
  assign mem[995] = 9'd7;
  assign mem[996] = 9'd6;
  assign mem[997] = 9'd5;
  assign mem[998] = 9'd4;
  assign mem[999] = 9'd3;
  assign mem[1000] = 9'd11;
  assign mem[1001] = 9'd10;
  assign mem[1002] = 9'd9;
  assign mem[1003] = 9'd8;
  assign mem[1004] = 9'd7;
  assign mem[1005] = 9'd6;
  assign mem[1006] = 9'd5;
  assign mem[1007] = 9'd4;
  assign mem[1008] = 9'd12;
  assign mem[1009] = 9'd11;
  assign mem[1010] = 9'd10;
  assign mem[1011] = 9'd9;
  assign mem[1012] = 9'd8;
  assign mem[1013] = 9'd7;
  assign mem[1014] = 9'd6;
  assign mem[1015] = 9'd5;
  assign mem[1016] = 9'd13;
  assign mem[1017] = 9'd12;
  assign mem[1018] = 9'd11;
  assign mem[1019] = 9'd10;
  assign mem[1020] = 9'd9;
  assign mem[1021] = 9'd8;
  assign mem[1022] = 9'd7;
  assign mem[1023] = 9'd6;
  assign mem[1024] = 9'd2;
  assign mem[1025] = 9'd3;
  assign mem[1026] = 9'd4;
  assign mem[1027] = 9'd5;
  assign mem[1028] = 9'd6;
  assign mem[1029] = 9'd7;
  assign mem[1030] = 9'd8;
  assign mem[1031] = 9'd9;
  assign mem[1032] = 9'd1;
  assign mem[1033] = 9'd2;
  assign mem[1034] = 9'd3;
  assign mem[1035] = 9'd4;
  assign mem[1036] = 9'd5;
  assign mem[1037] = 9'd6;
  assign mem[1038] = 9'd7;
  assign mem[1039] = 9'd8;
  assign mem[1040] = 9'd0;
  assign mem[1041] = 9'd1;
  assign mem[1042] = 9'd2;
  assign mem[1043] = 9'd3;
  assign mem[1044] = 9'd4;
  assign mem[1045] = 9'd5;
  assign mem[1046] = 9'd6;
  assign mem[1047] = 9'd7;
  assign mem[1048] = 9'd1;
  assign mem[1049] = 9'd2;
  assign mem[1050] = 9'd3;
  assign mem[1051] = 9'd4;
  assign mem[1052] = 9'd5;
  assign mem[1053] = 9'd6;
  assign mem[1054] = 9'd7;
  assign mem[1055] = 9'd8;
  assign mem[1056] = 9'd2;
  assign mem[1057] = 9'd3;
  assign mem[1058] = 9'd4;
  assign mem[1059] = 9'd5;
  assign mem[1060] = 9'd6;
  assign mem[1061] = 9'd7;
  assign mem[1062] = 9'd8;
  assign mem[1063] = 9'd9;
  assign mem[1064] = 9'd3;
  assign mem[1065] = 9'd4;
  assign mem[1066] = 9'd5;
  assign mem[1067] = 9'd6;
  assign mem[1068] = 9'd7;
  assign mem[1069] = 9'd8;
  assign mem[1070] = 9'd9;
  assign mem[1071] = 9'd10;
  assign mem[1072] = 9'd4;
  assign mem[1073] = 9'd5;
  assign mem[1074] = 9'd6;
  assign mem[1075] = 9'd7;
  assign mem[1076] = 9'd8;
  assign mem[1077] = 9'd9;
  assign mem[1078] = 9'd10;
  assign mem[1079] = 9'd11;
  assign mem[1080] = 9'd5;
  assign mem[1081] = 9'd6;
  assign mem[1082] = 9'd7;
  assign mem[1083] = 9'd8;
  assign mem[1084] = 9'd9;
  assign mem[1085] = 9'd10;
  assign mem[1086] = 9'd11;
  assign mem[1087] = 9'd12;
  assign mem[1088] = 9'd3;
  assign mem[1089] = 9'd2;
  assign mem[1090] = 9'd3;
  assign mem[1091] = 9'd4;
  assign mem[1092] = 9'd5;
  assign mem[1093] = 9'd6;
  assign mem[1094] = 9'd7;
  assign mem[1095] = 9'd8;
  assign mem[1096] = 9'd2;
  assign mem[1097] = 9'd1;
  assign mem[1098] = 9'd2;
  assign mem[1099] = 9'd3;
  assign mem[1100] = 9'd4;
  assign mem[1101] = 9'd5;
  assign mem[1102] = 9'd6;
  assign mem[1103] = 9'd7;
  assign mem[1104] = 9'd1;
  assign mem[1105] = 9'd0;
  assign mem[1106] = 9'd1;
  assign mem[1107] = 9'd2;
  assign mem[1108] = 9'd3;
  assign mem[1109] = 9'd4;
  assign mem[1110] = 9'd5;
  assign mem[1111] = 9'd6;
  assign mem[1112] = 9'd2;
  assign mem[1113] = 9'd1;
  assign mem[1114] = 9'd2;
  assign mem[1115] = 9'd3;
  assign mem[1116] = 9'd4;
  assign mem[1117] = 9'd5;
  assign mem[1118] = 9'd6;
  assign mem[1119] = 9'd7;
  assign mem[1120] = 9'd3;
  assign mem[1121] = 9'd2;
  assign mem[1122] = 9'd3;
  assign mem[1123] = 9'd4;
  assign mem[1124] = 9'd5;
  assign mem[1125] = 9'd6;
  assign mem[1126] = 9'd7;
  assign mem[1127] = 9'd8;
  assign mem[1128] = 9'd4;
  assign mem[1129] = 9'd3;
  assign mem[1130] = 9'd4;
  assign mem[1131] = 9'd5;
  assign mem[1132] = 9'd6;
  assign mem[1133] = 9'd7;
  assign mem[1134] = 9'd8;
  assign mem[1135] = 9'd9;
  assign mem[1136] = 9'd5;
  assign mem[1137] = 9'd4;
  assign mem[1138] = 9'd5;
  assign mem[1139] = 9'd6;
  assign mem[1140] = 9'd7;
  assign mem[1141] = 9'd8;
  assign mem[1142] = 9'd9;
  assign mem[1143] = 9'd10;
  assign mem[1144] = 9'd6;
  assign mem[1145] = 9'd5;
  assign mem[1146] = 9'd6;
  assign mem[1147] = 9'd7;
  assign mem[1148] = 9'd8;
  assign mem[1149] = 9'd9;
  assign mem[1150] = 9'd10;
  assign mem[1151] = 9'd11;
  assign mem[1152] = 9'd4;
  assign mem[1153] = 9'd3;
  assign mem[1154] = 9'd2;
  assign mem[1155] = 9'd3;
  assign mem[1156] = 9'd4;
  assign mem[1157] = 9'd5;
  assign mem[1158] = 9'd6;
  assign mem[1159] = 9'd7;
  assign mem[1160] = 9'd3;
  assign mem[1161] = 9'd2;
  assign mem[1162] = 9'd1;
  assign mem[1163] = 9'd2;
  assign mem[1164] = 9'd3;
  assign mem[1165] = 9'd4;
  assign mem[1166] = 9'd5;
  assign mem[1167] = 9'd6;
  assign mem[1168] = 9'd2;
  assign mem[1169] = 9'd1;
  assign mem[1170] = 9'd0;
  assign mem[1171] = 9'd1;
  assign mem[1172] = 9'd2;
  assign mem[1173] = 9'd3;
  assign mem[1174] = 9'd4;
  assign mem[1175] = 9'd5;
  assign mem[1176] = 9'd3;
  assign mem[1177] = 9'd2;
  assign mem[1178] = 9'd1;
  assign mem[1179] = 9'd2;
  assign mem[1180] = 9'd3;
  assign mem[1181] = 9'd4;
  assign mem[1182] = 9'd5;
  assign mem[1183] = 9'd6;
  assign mem[1184] = 9'd4;
  assign mem[1185] = 9'd3;
  assign mem[1186] = 9'd2;
  assign mem[1187] = 9'd3;
  assign mem[1188] = 9'd4;
  assign mem[1189] = 9'd5;
  assign mem[1190] = 9'd6;
  assign mem[1191] = 9'd7;
  assign mem[1192] = 9'd5;
  assign mem[1193] = 9'd4;
  assign mem[1194] = 9'd3;
  assign mem[1195] = 9'd4;
  assign mem[1196] = 9'd5;
  assign mem[1197] = 9'd6;
  assign mem[1198] = 9'd7;
  assign mem[1199] = 9'd8;
  assign mem[1200] = 9'd6;
  assign mem[1201] = 9'd5;
  assign mem[1202] = 9'd4;
  assign mem[1203] = 9'd5;
  assign mem[1204] = 9'd6;
  assign mem[1205] = 9'd7;
  assign mem[1206] = 9'd8;
  assign mem[1207] = 9'd9;
  assign mem[1208] = 9'd7;
  assign mem[1209] = 9'd6;
  assign mem[1210] = 9'd5;
  assign mem[1211] = 9'd6;
  assign mem[1212] = 9'd7;
  assign mem[1213] = 9'd8;
  assign mem[1214] = 9'd9;
  assign mem[1215] = 9'd10;
  assign mem[1216] = 9'd5;
  assign mem[1217] = 9'd4;
  assign mem[1218] = 9'd3;
  assign mem[1219] = 9'd2;
  assign mem[1220] = 9'd3;
  assign mem[1221] = 9'd4;
  assign mem[1222] = 9'd5;
  assign mem[1223] = 9'd6;
  assign mem[1224] = 9'd4;
  assign mem[1225] = 9'd3;
  assign mem[1226] = 9'd2;
  assign mem[1227] = 9'd1;
  assign mem[1228] = 9'd2;
  assign mem[1229] = 9'd3;
  assign mem[1230] = 9'd4;
  assign mem[1231] = 9'd5;
  assign mem[1232] = 9'd3;
  assign mem[1233] = 9'd2;
  assign mem[1234] = 9'd1;
  assign mem[1235] = 9'd0;
  assign mem[1236] = 9'd1;
  assign mem[1237] = 9'd2;
  assign mem[1238] = 9'd3;
  assign mem[1239] = 9'd4;
  assign mem[1240] = 9'd4;
  assign mem[1241] = 9'd3;
  assign mem[1242] = 9'd2;
  assign mem[1243] = 9'd1;
  assign mem[1244] = 9'd2;
  assign mem[1245] = 9'd3;
  assign mem[1246] = 9'd4;
  assign mem[1247] = 9'd5;
  assign mem[1248] = 9'd5;
  assign mem[1249] = 9'd4;
  assign mem[1250] = 9'd3;
  assign mem[1251] = 9'd2;
  assign mem[1252] = 9'd3;
  assign mem[1253] = 9'd4;
  assign mem[1254] = 9'd5;
  assign mem[1255] = 9'd6;
  assign mem[1256] = 9'd6;
  assign mem[1257] = 9'd5;
  assign mem[1258] = 9'd4;
  assign mem[1259] = 9'd3;
  assign mem[1260] = 9'd4;
  assign mem[1261] = 9'd5;
  assign mem[1262] = 9'd6;
  assign mem[1263] = 9'd7;
  assign mem[1264] = 9'd7;
  assign mem[1265] = 9'd6;
  assign mem[1266] = 9'd5;
  assign mem[1267] = 9'd4;
  assign mem[1268] = 9'd5;
  assign mem[1269] = 9'd6;
  assign mem[1270] = 9'd7;
  assign mem[1271] = 9'd8;
  assign mem[1272] = 9'd8;
  assign mem[1273] = 9'd7;
  assign mem[1274] = 9'd6;
  assign mem[1275] = 9'd5;
  assign mem[1276] = 9'd6;
  assign mem[1277] = 9'd7;
  assign mem[1278] = 9'd8;
  assign mem[1279] = 9'd9;
  assign mem[1280] = 9'd6;
  assign mem[1281] = 9'd5;
  assign mem[1282] = 9'd4;
  assign mem[1283] = 9'd3;
  assign mem[1284] = 9'd2;
  assign mem[1285] = 9'd3;
  assign mem[1286] = 9'd4;
  assign mem[1287] = 9'd5;
  assign mem[1288] = 9'd5;
  assign mem[1289] = 9'd4;
  assign mem[1290] = 9'd3;
  assign mem[1291] = 9'd2;
  assign mem[1292] = 9'd1;
  assign mem[1293] = 9'd2;
  assign mem[1294] = 9'd3;
  assign mem[1295] = 9'd4;
  assign mem[1296] = 9'd4;
  assign mem[1297] = 9'd3;
  assign mem[1298] = 9'd2;
  assign mem[1299] = 9'd1;
  assign mem[1300] = 9'd0;
  assign mem[1301] = 9'd1;
  assign mem[1302] = 9'd2;
  assign mem[1303] = 9'd3;
  assign mem[1304] = 9'd5;
  assign mem[1305] = 9'd4;
  assign mem[1306] = 9'd3;
  assign mem[1307] = 9'd2;
  assign mem[1308] = 9'd1;
  assign mem[1309] = 9'd2;
  assign mem[1310] = 9'd3;
  assign mem[1311] = 9'd4;
  assign mem[1312] = 9'd6;
  assign mem[1313] = 9'd5;
  assign mem[1314] = 9'd4;
  assign mem[1315] = 9'd3;
  assign mem[1316] = 9'd2;
  assign mem[1317] = 9'd3;
  assign mem[1318] = 9'd4;
  assign mem[1319] = 9'd5;
  assign mem[1320] = 9'd7;
  assign mem[1321] = 9'd6;
  assign mem[1322] = 9'd5;
  assign mem[1323] = 9'd4;
  assign mem[1324] = 9'd3;
  assign mem[1325] = 9'd4;
  assign mem[1326] = 9'd5;
  assign mem[1327] = 9'd6;
  assign mem[1328] = 9'd8;
  assign mem[1329] = 9'd7;
  assign mem[1330] = 9'd6;
  assign mem[1331] = 9'd5;
  assign mem[1332] = 9'd4;
  assign mem[1333] = 9'd5;
  assign mem[1334] = 9'd6;
  assign mem[1335] = 9'd7;
  assign mem[1336] = 9'd9;
  assign mem[1337] = 9'd8;
  assign mem[1338] = 9'd7;
  assign mem[1339] = 9'd6;
  assign mem[1340] = 9'd5;
  assign mem[1341] = 9'd6;
  assign mem[1342] = 9'd7;
  assign mem[1343] = 9'd8;
  assign mem[1344] = 9'd7;
  assign mem[1345] = 9'd6;
  assign mem[1346] = 9'd5;
  assign mem[1347] = 9'd4;
  assign mem[1348] = 9'd3;
  assign mem[1349] = 9'd2;
  assign mem[1350] = 9'd3;
  assign mem[1351] = 9'd4;
  assign mem[1352] = 9'd6;
  assign mem[1353] = 9'd5;
  assign mem[1354] = 9'd4;
  assign mem[1355] = 9'd3;
  assign mem[1356] = 9'd2;
  assign mem[1357] = 9'd1;
  assign mem[1358] = 9'd2;
  assign mem[1359] = 9'd3;
  assign mem[1360] = 9'd5;
  assign mem[1361] = 9'd4;
  assign mem[1362] = 9'd3;
  assign mem[1363] = 9'd2;
  assign mem[1364] = 9'd1;
  assign mem[1365] = 9'd0;
  assign mem[1366] = 9'd1;
  assign mem[1367] = 9'd2;
  assign mem[1368] = 9'd6;
  assign mem[1369] = 9'd5;
  assign mem[1370] = 9'd4;
  assign mem[1371] = 9'd3;
  assign mem[1372] = 9'd2;
  assign mem[1373] = 9'd1;
  assign mem[1374] = 9'd2;
  assign mem[1375] = 9'd3;
  assign mem[1376] = 9'd7;
  assign mem[1377] = 9'd6;
  assign mem[1378] = 9'd5;
  assign mem[1379] = 9'd4;
  assign mem[1380] = 9'd3;
  assign mem[1381] = 9'd2;
  assign mem[1382] = 9'd3;
  assign mem[1383] = 9'd4;
  assign mem[1384] = 9'd8;
  assign mem[1385] = 9'd7;
  assign mem[1386] = 9'd6;
  assign mem[1387] = 9'd5;
  assign mem[1388] = 9'd4;
  assign mem[1389] = 9'd3;
  assign mem[1390] = 9'd4;
  assign mem[1391] = 9'd5;
  assign mem[1392] = 9'd9;
  assign mem[1393] = 9'd8;
  assign mem[1394] = 9'd7;
  assign mem[1395] = 9'd6;
  assign mem[1396] = 9'd5;
  assign mem[1397] = 9'd4;
  assign mem[1398] = 9'd5;
  assign mem[1399] = 9'd6;
  assign mem[1400] = 9'd10;
  assign mem[1401] = 9'd9;
  assign mem[1402] = 9'd8;
  assign mem[1403] = 9'd7;
  assign mem[1404] = 9'd6;
  assign mem[1405] = 9'd5;
  assign mem[1406] = 9'd6;
  assign mem[1407] = 9'd7;
  assign mem[1408] = 9'd8;
  assign mem[1409] = 9'd7;
  assign mem[1410] = 9'd6;
  assign mem[1411] = 9'd5;
  assign mem[1412] = 9'd4;
  assign mem[1413] = 9'd3;
  assign mem[1414] = 9'd2;
  assign mem[1415] = 9'd3;
  assign mem[1416] = 9'd7;
  assign mem[1417] = 9'd6;
  assign mem[1418] = 9'd5;
  assign mem[1419] = 9'd4;
  assign mem[1420] = 9'd3;
  assign mem[1421] = 9'd2;
  assign mem[1422] = 9'd1;
  assign mem[1423] = 9'd2;
  assign mem[1424] = 9'd6;
  assign mem[1425] = 9'd5;
  assign mem[1426] = 9'd4;
  assign mem[1427] = 9'd3;
  assign mem[1428] = 9'd2;
  assign mem[1429] = 9'd1;
  assign mem[1430] = 9'd0;
  assign mem[1431] = 9'd1;
  assign mem[1432] = 9'd7;
  assign mem[1433] = 9'd6;
  assign mem[1434] = 9'd5;
  assign mem[1435] = 9'd4;
  assign mem[1436] = 9'd3;
  assign mem[1437] = 9'd2;
  assign mem[1438] = 9'd1;
  assign mem[1439] = 9'd2;
  assign mem[1440] = 9'd8;
  assign mem[1441] = 9'd7;
  assign mem[1442] = 9'd6;
  assign mem[1443] = 9'd5;
  assign mem[1444] = 9'd4;
  assign mem[1445] = 9'd3;
  assign mem[1446] = 9'd2;
  assign mem[1447] = 9'd3;
  assign mem[1448] = 9'd9;
  assign mem[1449] = 9'd8;
  assign mem[1450] = 9'd7;
  assign mem[1451] = 9'd6;
  assign mem[1452] = 9'd5;
  assign mem[1453] = 9'd4;
  assign mem[1454] = 9'd3;
  assign mem[1455] = 9'd4;
  assign mem[1456] = 9'd10;
  assign mem[1457] = 9'd9;
  assign mem[1458] = 9'd8;
  assign mem[1459] = 9'd7;
  assign mem[1460] = 9'd6;
  assign mem[1461] = 9'd5;
  assign mem[1462] = 9'd4;
  assign mem[1463] = 9'd5;
  assign mem[1464] = 9'd11;
  assign mem[1465] = 9'd10;
  assign mem[1466] = 9'd9;
  assign mem[1467] = 9'd8;
  assign mem[1468] = 9'd7;
  assign mem[1469] = 9'd6;
  assign mem[1470] = 9'd5;
  assign mem[1471] = 9'd6;
  assign mem[1472] = 9'd9;
  assign mem[1473] = 9'd8;
  assign mem[1474] = 9'd7;
  assign mem[1475] = 9'd6;
  assign mem[1476] = 9'd5;
  assign mem[1477] = 9'd4;
  assign mem[1478] = 9'd3;
  assign mem[1479] = 9'd2;
  assign mem[1480] = 9'd8;
  assign mem[1481] = 9'd7;
  assign mem[1482] = 9'd6;
  assign mem[1483] = 9'd5;
  assign mem[1484] = 9'd4;
  assign mem[1485] = 9'd3;
  assign mem[1486] = 9'd2;
  assign mem[1487] = 9'd1;
  assign mem[1488] = 9'd7;
  assign mem[1489] = 9'd6;
  assign mem[1490] = 9'd5;
  assign mem[1491] = 9'd4;
  assign mem[1492] = 9'd3;
  assign mem[1493] = 9'd2;
  assign mem[1494] = 9'd1;
  assign mem[1495] = 9'd0;
  assign mem[1496] = 9'd8;
  assign mem[1497] = 9'd7;
  assign mem[1498] = 9'd6;
  assign mem[1499] = 9'd5;
  assign mem[1500] = 9'd4;
  assign mem[1501] = 9'd3;
  assign mem[1502] = 9'd2;
  assign mem[1503] = 9'd1;
  assign mem[1504] = 9'd9;
  assign mem[1505] = 9'd8;
  assign mem[1506] = 9'd7;
  assign mem[1507] = 9'd6;
  assign mem[1508] = 9'd5;
  assign mem[1509] = 9'd4;
  assign mem[1510] = 9'd3;
  assign mem[1511] = 9'd2;
  assign mem[1512] = 9'd10;
  assign mem[1513] = 9'd9;
  assign mem[1514] = 9'd8;
  assign mem[1515] = 9'd7;
  assign mem[1516] = 9'd6;
  assign mem[1517] = 9'd5;
  assign mem[1518] = 9'd4;
  assign mem[1519] = 9'd3;
  assign mem[1520] = 9'd11;
  assign mem[1521] = 9'd10;
  assign mem[1522] = 9'd9;
  assign mem[1523] = 9'd8;
  assign mem[1524] = 9'd7;
  assign mem[1525] = 9'd6;
  assign mem[1526] = 9'd5;
  assign mem[1527] = 9'd4;
  assign mem[1528] = 9'd12;
  assign mem[1529] = 9'd11;
  assign mem[1530] = 9'd10;
  assign mem[1531] = 9'd9;
  assign mem[1532] = 9'd8;
  assign mem[1533] = 9'd7;
  assign mem[1534] = 9'd6;
  assign mem[1535] = 9'd5;
  assign mem[1536] = 9'd3;
  assign mem[1537] = 9'd4;
  assign mem[1538] = 9'd5;
  assign mem[1539] = 9'd6;
  assign mem[1540] = 9'd7;
  assign mem[1541] = 9'd8;
  assign mem[1542] = 9'd9;
  assign mem[1543] = 9'd10;
  assign mem[1544] = 9'd2;
  assign mem[1545] = 9'd3;
  assign mem[1546] = 9'd4;
  assign mem[1547] = 9'd5;
  assign mem[1548] = 9'd6;
  assign mem[1549] = 9'd7;
  assign mem[1550] = 9'd8;
  assign mem[1551] = 9'd9;
  assign mem[1552] = 9'd1;
  assign mem[1553] = 9'd2;
  assign mem[1554] = 9'd3;
  assign mem[1555] = 9'd4;
  assign mem[1556] = 9'd5;
  assign mem[1557] = 9'd6;
  assign mem[1558] = 9'd7;
  assign mem[1559] = 9'd8;
  assign mem[1560] = 9'd0;
  assign mem[1561] = 9'd1;
  assign mem[1562] = 9'd2;
  assign mem[1563] = 9'd3;
  assign mem[1564] = 9'd4;
  assign mem[1565] = 9'd5;
  assign mem[1566] = 9'd6;
  assign mem[1567] = 9'd7;
  assign mem[1568] = 9'd1;
  assign mem[1569] = 9'd2;
  assign mem[1570] = 9'd3;
  assign mem[1571] = 9'd4;
  assign mem[1572] = 9'd5;
  assign mem[1573] = 9'd6;
  assign mem[1574] = 9'd7;
  assign mem[1575] = 9'd8;
  assign mem[1576] = 9'd2;
  assign mem[1577] = 9'd3;
  assign mem[1578] = 9'd4;
  assign mem[1579] = 9'd5;
  assign mem[1580] = 9'd6;
  assign mem[1581] = 9'd7;
  assign mem[1582] = 9'd8;
  assign mem[1583] = 9'd9;
  assign mem[1584] = 9'd3;
  assign mem[1585] = 9'd4;
  assign mem[1586] = 9'd5;
  assign mem[1587] = 9'd6;
  assign mem[1588] = 9'd7;
  assign mem[1589] = 9'd8;
  assign mem[1590] = 9'd9;
  assign mem[1591] = 9'd10;
  assign mem[1592] = 9'd4;
  assign mem[1593] = 9'd5;
  assign mem[1594] = 9'd6;
  assign mem[1595] = 9'd7;
  assign mem[1596] = 9'd8;
  assign mem[1597] = 9'd9;
  assign mem[1598] = 9'd10;
  assign mem[1599] = 9'd11;
  assign mem[1600] = 9'd4;
  assign mem[1601] = 9'd3;
  assign mem[1602] = 9'd4;
  assign mem[1603] = 9'd5;
  assign mem[1604] = 9'd6;
  assign mem[1605] = 9'd7;
  assign mem[1606] = 9'd8;
  assign mem[1607] = 9'd9;
  assign mem[1608] = 9'd3;
  assign mem[1609] = 9'd2;
  assign mem[1610] = 9'd3;
  assign mem[1611] = 9'd4;
  assign mem[1612] = 9'd5;
  assign mem[1613] = 9'd6;
  assign mem[1614] = 9'd7;
  assign mem[1615] = 9'd8;
  assign mem[1616] = 9'd2;
  assign mem[1617] = 9'd1;
  assign mem[1618] = 9'd2;
  assign mem[1619] = 9'd3;
  assign mem[1620] = 9'd4;
  assign mem[1621] = 9'd5;
  assign mem[1622] = 9'd6;
  assign mem[1623] = 9'd7;
  assign mem[1624] = 9'd1;
  assign mem[1625] = 9'd0;
  assign mem[1626] = 9'd1;
  assign mem[1627] = 9'd2;
  assign mem[1628] = 9'd3;
  assign mem[1629] = 9'd4;
  assign mem[1630] = 9'd5;
  assign mem[1631] = 9'd6;
  assign mem[1632] = 9'd2;
  assign mem[1633] = 9'd1;
  assign mem[1634] = 9'd2;
  assign mem[1635] = 9'd3;
  assign mem[1636] = 9'd4;
  assign mem[1637] = 9'd5;
  assign mem[1638] = 9'd6;
  assign mem[1639] = 9'd7;
  assign mem[1640] = 9'd3;
  assign mem[1641] = 9'd2;
  assign mem[1642] = 9'd3;
  assign mem[1643] = 9'd4;
  assign mem[1644] = 9'd5;
  assign mem[1645] = 9'd6;
  assign mem[1646] = 9'd7;
  assign mem[1647] = 9'd8;
  assign mem[1648] = 9'd4;
  assign mem[1649] = 9'd3;
  assign mem[1650] = 9'd4;
  assign mem[1651] = 9'd5;
  assign mem[1652] = 9'd6;
  assign mem[1653] = 9'd7;
  assign mem[1654] = 9'd8;
  assign mem[1655] = 9'd9;
  assign mem[1656] = 9'd5;
  assign mem[1657] = 9'd4;
  assign mem[1658] = 9'd5;
  assign mem[1659] = 9'd6;
  assign mem[1660] = 9'd7;
  assign mem[1661] = 9'd8;
  assign mem[1662] = 9'd9;
  assign mem[1663] = 9'd10;
  assign mem[1664] = 9'd5;
  assign mem[1665] = 9'd4;
  assign mem[1666] = 9'd3;
  assign mem[1667] = 9'd4;
  assign mem[1668] = 9'd5;
  assign mem[1669] = 9'd6;
  assign mem[1670] = 9'd7;
  assign mem[1671] = 9'd8;
  assign mem[1672] = 9'd4;
  assign mem[1673] = 9'd3;
  assign mem[1674] = 9'd2;
  assign mem[1675] = 9'd3;
  assign mem[1676] = 9'd4;
  assign mem[1677] = 9'd5;
  assign mem[1678] = 9'd6;
  assign mem[1679] = 9'd7;
  assign mem[1680] = 9'd3;
  assign mem[1681] = 9'd2;
  assign mem[1682] = 9'd1;
  assign mem[1683] = 9'd2;
  assign mem[1684] = 9'd3;
  assign mem[1685] = 9'd4;
  assign mem[1686] = 9'd5;
  assign mem[1687] = 9'd6;
  assign mem[1688] = 9'd2;
  assign mem[1689] = 9'd1;
  assign mem[1690] = 9'd0;
  assign mem[1691] = 9'd1;
  assign mem[1692] = 9'd2;
  assign mem[1693] = 9'd3;
  assign mem[1694] = 9'd4;
  assign mem[1695] = 9'd5;
  assign mem[1696] = 9'd3;
  assign mem[1697] = 9'd2;
  assign mem[1698] = 9'd1;
  assign mem[1699] = 9'd2;
  assign mem[1700] = 9'd3;
  assign mem[1701] = 9'd4;
  assign mem[1702] = 9'd5;
  assign mem[1703] = 9'd6;
  assign mem[1704] = 9'd4;
  assign mem[1705] = 9'd3;
  assign mem[1706] = 9'd2;
  assign mem[1707] = 9'd3;
  assign mem[1708] = 9'd4;
  assign mem[1709] = 9'd5;
  assign mem[1710] = 9'd6;
  assign mem[1711] = 9'd7;
  assign mem[1712] = 9'd5;
  assign mem[1713] = 9'd4;
  assign mem[1714] = 9'd3;
  assign mem[1715] = 9'd4;
  assign mem[1716] = 9'd5;
  assign mem[1717] = 9'd6;
  assign mem[1718] = 9'd7;
  assign mem[1719] = 9'd8;
  assign mem[1720] = 9'd6;
  assign mem[1721] = 9'd5;
  assign mem[1722] = 9'd4;
  assign mem[1723] = 9'd5;
  assign mem[1724] = 9'd6;
  assign mem[1725] = 9'd7;
  assign mem[1726] = 9'd8;
  assign mem[1727] = 9'd9;
  assign mem[1728] = 9'd6;
  assign mem[1729] = 9'd5;
  assign mem[1730] = 9'd4;
  assign mem[1731] = 9'd3;
  assign mem[1732] = 9'd4;
  assign mem[1733] = 9'd5;
  assign mem[1734] = 9'd6;
  assign mem[1735] = 9'd7;
  assign mem[1736] = 9'd5;
  assign mem[1737] = 9'd4;
  assign mem[1738] = 9'd3;
  assign mem[1739] = 9'd2;
  assign mem[1740] = 9'd3;
  assign mem[1741] = 9'd4;
  assign mem[1742] = 9'd5;
  assign mem[1743] = 9'd6;
  assign mem[1744] = 9'd4;
  assign mem[1745] = 9'd3;
  assign mem[1746] = 9'd2;
  assign mem[1747] = 9'd1;
  assign mem[1748] = 9'd2;
  assign mem[1749] = 9'd3;
  assign mem[1750] = 9'd4;
  assign mem[1751] = 9'd5;
  assign mem[1752] = 9'd3;
  assign mem[1753] = 9'd2;
  assign mem[1754] = 9'd1;
  assign mem[1755] = 9'd0;
  assign mem[1756] = 9'd1;
  assign mem[1757] = 9'd2;
  assign mem[1758] = 9'd3;
  assign mem[1759] = 9'd4;
  assign mem[1760] = 9'd4;
  assign mem[1761] = 9'd3;
  assign mem[1762] = 9'd2;
  assign mem[1763] = 9'd1;
  assign mem[1764] = 9'd2;
  assign mem[1765] = 9'd3;
  assign mem[1766] = 9'd4;
  assign mem[1767] = 9'd5;
  assign mem[1768] = 9'd5;
  assign mem[1769] = 9'd4;
  assign mem[1770] = 9'd3;
  assign mem[1771] = 9'd2;
  assign mem[1772] = 9'd3;
  assign mem[1773] = 9'd4;
  assign mem[1774] = 9'd5;
  assign mem[1775] = 9'd6;
  assign mem[1776] = 9'd6;
  assign mem[1777] = 9'd5;
  assign mem[1778] = 9'd4;
  assign mem[1779] = 9'd3;
  assign mem[1780] = 9'd4;
  assign mem[1781] = 9'd5;
  assign mem[1782] = 9'd6;
  assign mem[1783] = 9'd7;
  assign mem[1784] = 9'd7;
  assign mem[1785] = 9'd6;
  assign mem[1786] = 9'd5;
  assign mem[1787] = 9'd4;
  assign mem[1788] = 9'd5;
  assign mem[1789] = 9'd6;
  assign mem[1790] = 9'd7;
  assign mem[1791] = 9'd8;
  assign mem[1792] = 9'd7;
  assign mem[1793] = 9'd6;
  assign mem[1794] = 9'd5;
  assign mem[1795] = 9'd4;
  assign mem[1796] = 9'd3;
  assign mem[1797] = 9'd4;
  assign mem[1798] = 9'd5;
  assign mem[1799] = 9'd6;
  assign mem[1800] = 9'd6;
  assign mem[1801] = 9'd5;
  assign mem[1802] = 9'd4;
  assign mem[1803] = 9'd3;
  assign mem[1804] = 9'd2;
  assign mem[1805] = 9'd3;
  assign mem[1806] = 9'd4;
  assign mem[1807] = 9'd5;
  assign mem[1808] = 9'd5;
  assign mem[1809] = 9'd4;
  assign mem[1810] = 9'd3;
  assign mem[1811] = 9'd2;
  assign mem[1812] = 9'd1;
  assign mem[1813] = 9'd2;
  assign mem[1814] = 9'd3;
  assign mem[1815] = 9'd4;
  assign mem[1816] = 9'd4;
  assign mem[1817] = 9'd3;
  assign mem[1818] = 9'd2;
  assign mem[1819] = 9'd1;
  assign mem[1820] = 9'd0;
  assign mem[1821] = 9'd1;
  assign mem[1822] = 9'd2;
  assign mem[1823] = 9'd3;
  assign mem[1824] = 9'd5;
  assign mem[1825] = 9'd4;
  assign mem[1826] = 9'd3;
  assign mem[1827] = 9'd2;
  assign mem[1828] = 9'd1;
  assign mem[1829] = 9'd2;
  assign mem[1830] = 9'd3;
  assign mem[1831] = 9'd4;
  assign mem[1832] = 9'd6;
  assign mem[1833] = 9'd5;
  assign mem[1834] = 9'd4;
  assign mem[1835] = 9'd3;
  assign mem[1836] = 9'd2;
  assign mem[1837] = 9'd3;
  assign mem[1838] = 9'd4;
  assign mem[1839] = 9'd5;
  assign mem[1840] = 9'd7;
  assign mem[1841] = 9'd6;
  assign mem[1842] = 9'd5;
  assign mem[1843] = 9'd4;
  assign mem[1844] = 9'd3;
  assign mem[1845] = 9'd4;
  assign mem[1846] = 9'd5;
  assign mem[1847] = 9'd6;
  assign mem[1848] = 9'd8;
  assign mem[1849] = 9'd7;
  assign mem[1850] = 9'd6;
  assign mem[1851] = 9'd5;
  assign mem[1852] = 9'd4;
  assign mem[1853] = 9'd5;
  assign mem[1854] = 9'd6;
  assign mem[1855] = 9'd7;
  assign mem[1856] = 9'd8;
  assign mem[1857] = 9'd7;
  assign mem[1858] = 9'd6;
  assign mem[1859] = 9'd5;
  assign mem[1860] = 9'd4;
  assign mem[1861] = 9'd3;
  assign mem[1862] = 9'd4;
  assign mem[1863] = 9'd5;
  assign mem[1864] = 9'd7;
  assign mem[1865] = 9'd6;
  assign mem[1866] = 9'd5;
  assign mem[1867] = 9'd4;
  assign mem[1868] = 9'd3;
  assign mem[1869] = 9'd2;
  assign mem[1870] = 9'd3;
  assign mem[1871] = 9'd4;
  assign mem[1872] = 9'd6;
  assign mem[1873] = 9'd5;
  assign mem[1874] = 9'd4;
  assign mem[1875] = 9'd3;
  assign mem[1876] = 9'd2;
  assign mem[1877] = 9'd1;
  assign mem[1878] = 9'd2;
  assign mem[1879] = 9'd3;
  assign mem[1880] = 9'd5;
  assign mem[1881] = 9'd4;
  assign mem[1882] = 9'd3;
  assign mem[1883] = 9'd2;
  assign mem[1884] = 9'd1;
  assign mem[1885] = 9'd0;
  assign mem[1886] = 9'd1;
  assign mem[1887] = 9'd2;
  assign mem[1888] = 9'd6;
  assign mem[1889] = 9'd5;
  assign mem[1890] = 9'd4;
  assign mem[1891] = 9'd3;
  assign mem[1892] = 9'd2;
  assign mem[1893] = 9'd1;
  assign mem[1894] = 9'd2;
  assign mem[1895] = 9'd3;
  assign mem[1896] = 9'd7;
  assign mem[1897] = 9'd6;
  assign mem[1898] = 9'd5;
  assign mem[1899] = 9'd4;
  assign mem[1900] = 9'd3;
  assign mem[1901] = 9'd2;
  assign mem[1902] = 9'd3;
  assign mem[1903] = 9'd4;
  assign mem[1904] = 9'd8;
  assign mem[1905] = 9'd7;
  assign mem[1906] = 9'd6;
  assign mem[1907] = 9'd5;
  assign mem[1908] = 9'd4;
  assign mem[1909] = 9'd3;
  assign mem[1910] = 9'd4;
  assign mem[1911] = 9'd5;
  assign mem[1912] = 9'd9;
  assign mem[1913] = 9'd8;
  assign mem[1914] = 9'd7;
  assign mem[1915] = 9'd6;
  assign mem[1916] = 9'd5;
  assign mem[1917] = 9'd4;
  assign mem[1918] = 9'd5;
  assign mem[1919] = 9'd6;
  assign mem[1920] = 9'd9;
  assign mem[1921] = 9'd8;
  assign mem[1922] = 9'd7;
  assign mem[1923] = 9'd6;
  assign mem[1924] = 9'd5;
  assign mem[1925] = 9'd4;
  assign mem[1926] = 9'd3;
  assign mem[1927] = 9'd4;
  assign mem[1928] = 9'd8;
  assign mem[1929] = 9'd7;
  assign mem[1930] = 9'd6;
  assign mem[1931] = 9'd5;
  assign mem[1932] = 9'd4;
  assign mem[1933] = 9'd3;
  assign mem[1934] = 9'd2;
  assign mem[1935] = 9'd3;
  assign mem[1936] = 9'd7;
  assign mem[1937] = 9'd6;
  assign mem[1938] = 9'd5;
  assign mem[1939] = 9'd4;
  assign mem[1940] = 9'd3;
  assign mem[1941] = 9'd2;
  assign mem[1942] = 9'd1;
  assign mem[1943] = 9'd2;
  assign mem[1944] = 9'd6;
  assign mem[1945] = 9'd5;
  assign mem[1946] = 9'd4;
  assign mem[1947] = 9'd3;
  assign mem[1948] = 9'd2;
  assign mem[1949] = 9'd1;
  assign mem[1950] = 9'd0;
  assign mem[1951] = 9'd1;
  assign mem[1952] = 9'd7;
  assign mem[1953] = 9'd6;
  assign mem[1954] = 9'd5;
  assign mem[1955] = 9'd4;
  assign mem[1956] = 9'd3;
  assign mem[1957] = 9'd2;
  assign mem[1958] = 9'd1;
  assign mem[1959] = 9'd2;
  assign mem[1960] = 9'd8;
  assign mem[1961] = 9'd7;
  assign mem[1962] = 9'd6;
  assign mem[1963] = 9'd5;
  assign mem[1964] = 9'd4;
  assign mem[1965] = 9'd3;
  assign mem[1966] = 9'd2;
  assign mem[1967] = 9'd3;
  assign mem[1968] = 9'd9;
  assign mem[1969] = 9'd8;
  assign mem[1970] = 9'd7;
  assign mem[1971] = 9'd6;
  assign mem[1972] = 9'd5;
  assign mem[1973] = 9'd4;
  assign mem[1974] = 9'd3;
  assign mem[1975] = 9'd4;
  assign mem[1976] = 9'd10;
  assign mem[1977] = 9'd9;
  assign mem[1978] = 9'd8;
  assign mem[1979] = 9'd7;
  assign mem[1980] = 9'd6;
  assign mem[1981] = 9'd5;
  assign mem[1982] = 9'd4;
  assign mem[1983] = 9'd5;
  assign mem[1984] = 9'd10;
  assign mem[1985] = 9'd9;
  assign mem[1986] = 9'd8;
  assign mem[1987] = 9'd7;
  assign mem[1988] = 9'd6;
  assign mem[1989] = 9'd5;
  assign mem[1990] = 9'd4;
  assign mem[1991] = 9'd3;
  assign mem[1992] = 9'd9;
  assign mem[1993] = 9'd8;
  assign mem[1994] = 9'd7;
  assign mem[1995] = 9'd6;
  assign mem[1996] = 9'd5;
  assign mem[1997] = 9'd4;
  assign mem[1998] = 9'd3;
  assign mem[1999] = 9'd2;
  assign mem[2000] = 9'd8;
  assign mem[2001] = 9'd7;
  assign mem[2002] = 9'd6;
  assign mem[2003] = 9'd5;
  assign mem[2004] = 9'd4;
  assign mem[2005] = 9'd3;
  assign mem[2006] = 9'd2;
  assign mem[2007] = 9'd1;
  assign mem[2008] = 9'd7;
  assign mem[2009] = 9'd6;
  assign mem[2010] = 9'd5;
  assign mem[2011] = 9'd4;
  assign mem[2012] = 9'd3;
  assign mem[2013] = 9'd2;
  assign mem[2014] = 9'd1;
  assign mem[2015] = 9'd0;
  assign mem[2016] = 9'd8;
  assign mem[2017] = 9'd7;
  assign mem[2018] = 9'd6;
  assign mem[2019] = 9'd5;
  assign mem[2020] = 9'd4;
  assign mem[2021] = 9'd3;
  assign mem[2022] = 9'd2;
  assign mem[2023] = 9'd1;
  assign mem[2024] = 9'd9;
  assign mem[2025] = 9'd8;
  assign mem[2026] = 9'd7;
  assign mem[2027] = 9'd6;
  assign mem[2028] = 9'd5;
  assign mem[2029] = 9'd4;
  assign mem[2030] = 9'd3;
  assign mem[2031] = 9'd2;
  assign mem[2032] = 9'd10;
  assign mem[2033] = 9'd9;
  assign mem[2034] = 9'd8;
  assign mem[2035] = 9'd7;
  assign mem[2036] = 9'd6;
  assign mem[2037] = 9'd5;
  assign mem[2038] = 9'd4;
  assign mem[2039] = 9'd3;
  assign mem[2040] = 9'd11;
  assign mem[2041] = 9'd10;
  assign mem[2042] = 9'd9;
  assign mem[2043] = 9'd8;
  assign mem[2044] = 9'd7;
  assign mem[2045] = 9'd6;
  assign mem[2046] = 9'd5;
  assign mem[2047] = 9'd4;
  assign mem[2048] = 9'd4;
  assign mem[2049] = 9'd5;
  assign mem[2050] = 9'd6;
  assign mem[2051] = 9'd7;
  assign mem[2052] = 9'd8;
  assign mem[2053] = 9'd9;
  assign mem[2054] = 9'd10;
  assign mem[2055] = 9'd11;
  assign mem[2056] = 9'd3;
  assign mem[2057] = 9'd4;
  assign mem[2058] = 9'd5;
  assign mem[2059] = 9'd6;
  assign mem[2060] = 9'd7;
  assign mem[2061] = 9'd8;
  assign mem[2062] = 9'd9;
  assign mem[2063] = 9'd10;
  assign mem[2064] = 9'd2;
  assign mem[2065] = 9'd3;
  assign mem[2066] = 9'd4;
  assign mem[2067] = 9'd5;
  assign mem[2068] = 9'd6;
  assign mem[2069] = 9'd7;
  assign mem[2070] = 9'd8;
  assign mem[2071] = 9'd9;
  assign mem[2072] = 9'd1;
  assign mem[2073] = 9'd2;
  assign mem[2074] = 9'd3;
  assign mem[2075] = 9'd4;
  assign mem[2076] = 9'd5;
  assign mem[2077] = 9'd6;
  assign mem[2078] = 9'd7;
  assign mem[2079] = 9'd8;
  assign mem[2080] = 9'd0;
  assign mem[2081] = 9'd1;
  assign mem[2082] = 9'd2;
  assign mem[2083] = 9'd3;
  assign mem[2084] = 9'd4;
  assign mem[2085] = 9'd5;
  assign mem[2086] = 9'd6;
  assign mem[2087] = 9'd7;
  assign mem[2088] = 9'd1;
  assign mem[2089] = 9'd2;
  assign mem[2090] = 9'd3;
  assign mem[2091] = 9'd4;
  assign mem[2092] = 9'd5;
  assign mem[2093] = 9'd6;
  assign mem[2094] = 9'd7;
  assign mem[2095] = 9'd8;
  assign mem[2096] = 9'd2;
  assign mem[2097] = 9'd3;
  assign mem[2098] = 9'd4;
  assign mem[2099] = 9'd5;
  assign mem[2100] = 9'd6;
  assign mem[2101] = 9'd7;
  assign mem[2102] = 9'd8;
  assign mem[2103] = 9'd9;
  assign mem[2104] = 9'd3;
  assign mem[2105] = 9'd4;
  assign mem[2106] = 9'd5;
  assign mem[2107] = 9'd6;
  assign mem[2108] = 9'd7;
  assign mem[2109] = 9'd8;
  assign mem[2110] = 9'd9;
  assign mem[2111] = 9'd10;
  assign mem[2112] = 9'd5;
  assign mem[2113] = 9'd4;
  assign mem[2114] = 9'd5;
  assign mem[2115] = 9'd6;
  assign mem[2116] = 9'd7;
  assign mem[2117] = 9'd8;
  assign mem[2118] = 9'd9;
  assign mem[2119] = 9'd10;
  assign mem[2120] = 9'd4;
  assign mem[2121] = 9'd3;
  assign mem[2122] = 9'd4;
  assign mem[2123] = 9'd5;
  assign mem[2124] = 9'd6;
  assign mem[2125] = 9'd7;
  assign mem[2126] = 9'd8;
  assign mem[2127] = 9'd9;
  assign mem[2128] = 9'd3;
  assign mem[2129] = 9'd2;
  assign mem[2130] = 9'd3;
  assign mem[2131] = 9'd4;
  assign mem[2132] = 9'd5;
  assign mem[2133] = 9'd6;
  assign mem[2134] = 9'd7;
  assign mem[2135] = 9'd8;
  assign mem[2136] = 9'd2;
  assign mem[2137] = 9'd1;
  assign mem[2138] = 9'd2;
  assign mem[2139] = 9'd3;
  assign mem[2140] = 9'd4;
  assign mem[2141] = 9'd5;
  assign mem[2142] = 9'd6;
  assign mem[2143] = 9'd7;
  assign mem[2144] = 9'd1;
  assign mem[2145] = 9'd0;
  assign mem[2146] = 9'd1;
  assign mem[2147] = 9'd2;
  assign mem[2148] = 9'd3;
  assign mem[2149] = 9'd4;
  assign mem[2150] = 9'd5;
  assign mem[2151] = 9'd6;
  assign mem[2152] = 9'd2;
  assign mem[2153] = 9'd1;
  assign mem[2154] = 9'd2;
  assign mem[2155] = 9'd3;
  assign mem[2156] = 9'd4;
  assign mem[2157] = 9'd5;
  assign mem[2158] = 9'd6;
  assign mem[2159] = 9'd7;
  assign mem[2160] = 9'd3;
  assign mem[2161] = 9'd2;
  assign mem[2162] = 9'd3;
  assign mem[2163] = 9'd4;
  assign mem[2164] = 9'd5;
  assign mem[2165] = 9'd6;
  assign mem[2166] = 9'd7;
  assign mem[2167] = 9'd8;
  assign mem[2168] = 9'd4;
  assign mem[2169] = 9'd3;
  assign mem[2170] = 9'd4;
  assign mem[2171] = 9'd5;
  assign mem[2172] = 9'd6;
  assign mem[2173] = 9'd7;
  assign mem[2174] = 9'd8;
  assign mem[2175] = 9'd9;
  assign mem[2176] = 9'd6;
  assign mem[2177] = 9'd5;
  assign mem[2178] = 9'd4;
  assign mem[2179] = 9'd5;
  assign mem[2180] = 9'd6;
  assign mem[2181] = 9'd7;
  assign mem[2182] = 9'd8;
  assign mem[2183] = 9'd9;
  assign mem[2184] = 9'd5;
  assign mem[2185] = 9'd4;
  assign mem[2186] = 9'd3;
  assign mem[2187] = 9'd4;
  assign mem[2188] = 9'd5;
  assign mem[2189] = 9'd6;
  assign mem[2190] = 9'd7;
  assign mem[2191] = 9'd8;
  assign mem[2192] = 9'd4;
  assign mem[2193] = 9'd3;
  assign mem[2194] = 9'd2;
  assign mem[2195] = 9'd3;
  assign mem[2196] = 9'd4;
  assign mem[2197] = 9'd5;
  assign mem[2198] = 9'd6;
  assign mem[2199] = 9'd7;
  assign mem[2200] = 9'd3;
  assign mem[2201] = 9'd2;
  assign mem[2202] = 9'd1;
  assign mem[2203] = 9'd2;
  assign mem[2204] = 9'd3;
  assign mem[2205] = 9'd4;
  assign mem[2206] = 9'd5;
  assign mem[2207] = 9'd6;
  assign mem[2208] = 9'd2;
  assign mem[2209] = 9'd1;
  assign mem[2210] = 9'd0;
  assign mem[2211] = 9'd1;
  assign mem[2212] = 9'd2;
  assign mem[2213] = 9'd3;
  assign mem[2214] = 9'd4;
  assign mem[2215] = 9'd5;
  assign mem[2216] = 9'd3;
  assign mem[2217] = 9'd2;
  assign mem[2218] = 9'd1;
  assign mem[2219] = 9'd2;
  assign mem[2220] = 9'd3;
  assign mem[2221] = 9'd4;
  assign mem[2222] = 9'd5;
  assign mem[2223] = 9'd6;
  assign mem[2224] = 9'd4;
  assign mem[2225] = 9'd3;
  assign mem[2226] = 9'd2;
  assign mem[2227] = 9'd3;
  assign mem[2228] = 9'd4;
  assign mem[2229] = 9'd5;
  assign mem[2230] = 9'd6;
  assign mem[2231] = 9'd7;
  assign mem[2232] = 9'd5;
  assign mem[2233] = 9'd4;
  assign mem[2234] = 9'd3;
  assign mem[2235] = 9'd4;
  assign mem[2236] = 9'd5;
  assign mem[2237] = 9'd6;
  assign mem[2238] = 9'd7;
  assign mem[2239] = 9'd8;
  assign mem[2240] = 9'd7;
  assign mem[2241] = 9'd6;
  assign mem[2242] = 9'd5;
  assign mem[2243] = 9'd4;
  assign mem[2244] = 9'd5;
  assign mem[2245] = 9'd6;
  assign mem[2246] = 9'd7;
  assign mem[2247] = 9'd8;
  assign mem[2248] = 9'd6;
  assign mem[2249] = 9'd5;
  assign mem[2250] = 9'd4;
  assign mem[2251] = 9'd3;
  assign mem[2252] = 9'd4;
  assign mem[2253] = 9'd5;
  assign mem[2254] = 9'd6;
  assign mem[2255] = 9'd7;
  assign mem[2256] = 9'd5;
  assign mem[2257] = 9'd4;
  assign mem[2258] = 9'd3;
  assign mem[2259] = 9'd2;
  assign mem[2260] = 9'd3;
  assign mem[2261] = 9'd4;
  assign mem[2262] = 9'd5;
  assign mem[2263] = 9'd6;
  assign mem[2264] = 9'd4;
  assign mem[2265] = 9'd3;
  assign mem[2266] = 9'd2;
  assign mem[2267] = 9'd1;
  assign mem[2268] = 9'd2;
  assign mem[2269] = 9'd3;
  assign mem[2270] = 9'd4;
  assign mem[2271] = 9'd5;
  assign mem[2272] = 9'd3;
  assign mem[2273] = 9'd2;
  assign mem[2274] = 9'd1;
  assign mem[2275] = 9'd0;
  assign mem[2276] = 9'd1;
  assign mem[2277] = 9'd2;
  assign mem[2278] = 9'd3;
  assign mem[2279] = 9'd4;
  assign mem[2280] = 9'd4;
  assign mem[2281] = 9'd3;
  assign mem[2282] = 9'd2;
  assign mem[2283] = 9'd1;
  assign mem[2284] = 9'd2;
  assign mem[2285] = 9'd3;
  assign mem[2286] = 9'd4;
  assign mem[2287] = 9'd5;
  assign mem[2288] = 9'd5;
  assign mem[2289] = 9'd4;
  assign mem[2290] = 9'd3;
  assign mem[2291] = 9'd2;
  assign mem[2292] = 9'd3;
  assign mem[2293] = 9'd4;
  assign mem[2294] = 9'd5;
  assign mem[2295] = 9'd6;
  assign mem[2296] = 9'd6;
  assign mem[2297] = 9'd5;
  assign mem[2298] = 9'd4;
  assign mem[2299] = 9'd3;
  assign mem[2300] = 9'd4;
  assign mem[2301] = 9'd5;
  assign mem[2302] = 9'd6;
  assign mem[2303] = 9'd7;
  assign mem[2304] = 9'd8;
  assign mem[2305] = 9'd7;
  assign mem[2306] = 9'd6;
  assign mem[2307] = 9'd5;
  assign mem[2308] = 9'd4;
  assign mem[2309] = 9'd5;
  assign mem[2310] = 9'd6;
  assign mem[2311] = 9'd7;
  assign mem[2312] = 9'd7;
  assign mem[2313] = 9'd6;
  assign mem[2314] = 9'd5;
  assign mem[2315] = 9'd4;
  assign mem[2316] = 9'd3;
  assign mem[2317] = 9'd4;
  assign mem[2318] = 9'd5;
  assign mem[2319] = 9'd6;
  assign mem[2320] = 9'd6;
  assign mem[2321] = 9'd5;
  assign mem[2322] = 9'd4;
  assign mem[2323] = 9'd3;
  assign mem[2324] = 9'd2;
  assign mem[2325] = 9'd3;
  assign mem[2326] = 9'd4;
  assign mem[2327] = 9'd5;
  assign mem[2328] = 9'd5;
  assign mem[2329] = 9'd4;
  assign mem[2330] = 9'd3;
  assign mem[2331] = 9'd2;
  assign mem[2332] = 9'd1;
  assign mem[2333] = 9'd2;
  assign mem[2334] = 9'd3;
  assign mem[2335] = 9'd4;
  assign mem[2336] = 9'd4;
  assign mem[2337] = 9'd3;
  assign mem[2338] = 9'd2;
  assign mem[2339] = 9'd1;
  assign mem[2340] = 9'd0;
  assign mem[2341] = 9'd1;
  assign mem[2342] = 9'd2;
  assign mem[2343] = 9'd3;
  assign mem[2344] = 9'd5;
  assign mem[2345] = 9'd4;
  assign mem[2346] = 9'd3;
  assign mem[2347] = 9'd2;
  assign mem[2348] = 9'd1;
  assign mem[2349] = 9'd2;
  assign mem[2350] = 9'd3;
  assign mem[2351] = 9'd4;
  assign mem[2352] = 9'd6;
  assign mem[2353] = 9'd5;
  assign mem[2354] = 9'd4;
  assign mem[2355] = 9'd3;
  assign mem[2356] = 9'd2;
  assign mem[2357] = 9'd3;
  assign mem[2358] = 9'd4;
  assign mem[2359] = 9'd5;
  assign mem[2360] = 9'd7;
  assign mem[2361] = 9'd6;
  assign mem[2362] = 9'd5;
  assign mem[2363] = 9'd4;
  assign mem[2364] = 9'd3;
  assign mem[2365] = 9'd4;
  assign mem[2366] = 9'd5;
  assign mem[2367] = 9'd6;
  assign mem[2368] = 9'd9;
  assign mem[2369] = 9'd8;
  assign mem[2370] = 9'd7;
  assign mem[2371] = 9'd6;
  assign mem[2372] = 9'd5;
  assign mem[2373] = 9'd4;
  assign mem[2374] = 9'd5;
  assign mem[2375] = 9'd6;
  assign mem[2376] = 9'd8;
  assign mem[2377] = 9'd7;
  assign mem[2378] = 9'd6;
  assign mem[2379] = 9'd5;
  assign mem[2380] = 9'd4;
  assign mem[2381] = 9'd3;
  assign mem[2382] = 9'd4;
  assign mem[2383] = 9'd5;
  assign mem[2384] = 9'd7;
  assign mem[2385] = 9'd6;
  assign mem[2386] = 9'd5;
  assign mem[2387] = 9'd4;
  assign mem[2388] = 9'd3;
  assign mem[2389] = 9'd2;
  assign mem[2390] = 9'd3;
  assign mem[2391] = 9'd4;
  assign mem[2392] = 9'd6;
  assign mem[2393] = 9'd5;
  assign mem[2394] = 9'd4;
  assign mem[2395] = 9'd3;
  assign mem[2396] = 9'd2;
  assign mem[2397] = 9'd1;
  assign mem[2398] = 9'd2;
  assign mem[2399] = 9'd3;
  assign mem[2400] = 9'd5;
  assign mem[2401] = 9'd4;
  assign mem[2402] = 9'd3;
  assign mem[2403] = 9'd2;
  assign mem[2404] = 9'd1;
  assign mem[2405] = 9'd0;
  assign mem[2406] = 9'd1;
  assign mem[2407] = 9'd2;
  assign mem[2408] = 9'd6;
  assign mem[2409] = 9'd5;
  assign mem[2410] = 9'd4;
  assign mem[2411] = 9'd3;
  assign mem[2412] = 9'd2;
  assign mem[2413] = 9'd1;
  assign mem[2414] = 9'd2;
  assign mem[2415] = 9'd3;
  assign mem[2416] = 9'd7;
  assign mem[2417] = 9'd6;
  assign mem[2418] = 9'd5;
  assign mem[2419] = 9'd4;
  assign mem[2420] = 9'd3;
  assign mem[2421] = 9'd2;
  assign mem[2422] = 9'd3;
  assign mem[2423] = 9'd4;
  assign mem[2424] = 9'd8;
  assign mem[2425] = 9'd7;
  assign mem[2426] = 9'd6;
  assign mem[2427] = 9'd5;
  assign mem[2428] = 9'd4;
  assign mem[2429] = 9'd3;
  assign mem[2430] = 9'd4;
  assign mem[2431] = 9'd5;
  assign mem[2432] = 9'd10;
  assign mem[2433] = 9'd9;
  assign mem[2434] = 9'd8;
  assign mem[2435] = 9'd7;
  assign mem[2436] = 9'd6;
  assign mem[2437] = 9'd5;
  assign mem[2438] = 9'd4;
  assign mem[2439] = 9'd5;
  assign mem[2440] = 9'd9;
  assign mem[2441] = 9'd8;
  assign mem[2442] = 9'd7;
  assign mem[2443] = 9'd6;
  assign mem[2444] = 9'd5;
  assign mem[2445] = 9'd4;
  assign mem[2446] = 9'd3;
  assign mem[2447] = 9'd4;
  assign mem[2448] = 9'd8;
  assign mem[2449] = 9'd7;
  assign mem[2450] = 9'd6;
  assign mem[2451] = 9'd5;
  assign mem[2452] = 9'd4;
  assign mem[2453] = 9'd3;
  assign mem[2454] = 9'd2;
  assign mem[2455] = 9'd3;
  assign mem[2456] = 9'd7;
  assign mem[2457] = 9'd6;
  assign mem[2458] = 9'd5;
  assign mem[2459] = 9'd4;
  assign mem[2460] = 9'd3;
  assign mem[2461] = 9'd2;
  assign mem[2462] = 9'd1;
  assign mem[2463] = 9'd2;
  assign mem[2464] = 9'd6;
  assign mem[2465] = 9'd5;
  assign mem[2466] = 9'd4;
  assign mem[2467] = 9'd3;
  assign mem[2468] = 9'd2;
  assign mem[2469] = 9'd1;
  assign mem[2470] = 9'd0;
  assign mem[2471] = 9'd1;
  assign mem[2472] = 9'd7;
  assign mem[2473] = 9'd6;
  assign mem[2474] = 9'd5;
  assign mem[2475] = 9'd4;
  assign mem[2476] = 9'd3;
  assign mem[2477] = 9'd2;
  assign mem[2478] = 9'd1;
  assign mem[2479] = 9'd2;
  assign mem[2480] = 9'd8;
  assign mem[2481] = 9'd7;
  assign mem[2482] = 9'd6;
  assign mem[2483] = 9'd5;
  assign mem[2484] = 9'd4;
  assign mem[2485] = 9'd3;
  assign mem[2486] = 9'd2;
  assign mem[2487] = 9'd3;
  assign mem[2488] = 9'd9;
  assign mem[2489] = 9'd8;
  assign mem[2490] = 9'd7;
  assign mem[2491] = 9'd6;
  assign mem[2492] = 9'd5;
  assign mem[2493] = 9'd4;
  assign mem[2494] = 9'd3;
  assign mem[2495] = 9'd4;
  assign mem[2496] = 9'd11;
  assign mem[2497] = 9'd10;
  assign mem[2498] = 9'd9;
  assign mem[2499] = 9'd8;
  assign mem[2500] = 9'd7;
  assign mem[2501] = 9'd6;
  assign mem[2502] = 9'd5;
  assign mem[2503] = 9'd4;
  assign mem[2504] = 9'd10;
  assign mem[2505] = 9'd9;
  assign mem[2506] = 9'd8;
  assign mem[2507] = 9'd7;
  assign mem[2508] = 9'd6;
  assign mem[2509] = 9'd5;
  assign mem[2510] = 9'd4;
  assign mem[2511] = 9'd3;
  assign mem[2512] = 9'd9;
  assign mem[2513] = 9'd8;
  assign mem[2514] = 9'd7;
  assign mem[2515] = 9'd6;
  assign mem[2516] = 9'd5;
  assign mem[2517] = 9'd4;
  assign mem[2518] = 9'd3;
  assign mem[2519] = 9'd2;
  assign mem[2520] = 9'd8;
  assign mem[2521] = 9'd7;
  assign mem[2522] = 9'd6;
  assign mem[2523] = 9'd5;
  assign mem[2524] = 9'd4;
  assign mem[2525] = 9'd3;
  assign mem[2526] = 9'd2;
  assign mem[2527] = 9'd1;
  assign mem[2528] = 9'd7;
  assign mem[2529] = 9'd6;
  assign mem[2530] = 9'd5;
  assign mem[2531] = 9'd4;
  assign mem[2532] = 9'd3;
  assign mem[2533] = 9'd2;
  assign mem[2534] = 9'd1;
  assign mem[2535] = 9'd0;
  assign mem[2536] = 9'd8;
  assign mem[2537] = 9'd7;
  assign mem[2538] = 9'd6;
  assign mem[2539] = 9'd5;
  assign mem[2540] = 9'd4;
  assign mem[2541] = 9'd3;
  assign mem[2542] = 9'd2;
  assign mem[2543] = 9'd1;
  assign mem[2544] = 9'd9;
  assign mem[2545] = 9'd8;
  assign mem[2546] = 9'd7;
  assign mem[2547] = 9'd6;
  assign mem[2548] = 9'd5;
  assign mem[2549] = 9'd4;
  assign mem[2550] = 9'd3;
  assign mem[2551] = 9'd2;
  assign mem[2552] = 9'd10;
  assign mem[2553] = 9'd9;
  assign mem[2554] = 9'd8;
  assign mem[2555] = 9'd7;
  assign mem[2556] = 9'd6;
  assign mem[2557] = 9'd5;
  assign mem[2558] = 9'd4;
  assign mem[2559] = 9'd3;
  assign mem[2560] = 9'd5;
  assign mem[2561] = 9'd6;
  assign mem[2562] = 9'd7;
  assign mem[2563] = 9'd8;
  assign mem[2564] = 9'd9;
  assign mem[2565] = 9'd10;
  assign mem[2566] = 9'd11;
  assign mem[2567] = 9'd12;
  assign mem[2568] = 9'd4;
  assign mem[2569] = 9'd5;
  assign mem[2570] = 9'd6;
  assign mem[2571] = 9'd7;
  assign mem[2572] = 9'd8;
  assign mem[2573] = 9'd9;
  assign mem[2574] = 9'd10;
  assign mem[2575] = 9'd11;
  assign mem[2576] = 9'd3;
  assign mem[2577] = 9'd4;
  assign mem[2578] = 9'd5;
  assign mem[2579] = 9'd6;
  assign mem[2580] = 9'd7;
  assign mem[2581] = 9'd8;
  assign mem[2582] = 9'd9;
  assign mem[2583] = 9'd10;
  assign mem[2584] = 9'd2;
  assign mem[2585] = 9'd3;
  assign mem[2586] = 9'd4;
  assign mem[2587] = 9'd5;
  assign mem[2588] = 9'd6;
  assign mem[2589] = 9'd7;
  assign mem[2590] = 9'd8;
  assign mem[2591] = 9'd9;
  assign mem[2592] = 9'd1;
  assign mem[2593] = 9'd2;
  assign mem[2594] = 9'd3;
  assign mem[2595] = 9'd4;
  assign mem[2596] = 9'd5;
  assign mem[2597] = 9'd6;
  assign mem[2598] = 9'd7;
  assign mem[2599] = 9'd8;
  assign mem[2600] = 9'd0;
  assign mem[2601] = 9'd1;
  assign mem[2602] = 9'd2;
  assign mem[2603] = 9'd3;
  assign mem[2604] = 9'd4;
  assign mem[2605] = 9'd5;
  assign mem[2606] = 9'd6;
  assign mem[2607] = 9'd7;
  assign mem[2608] = 9'd1;
  assign mem[2609] = 9'd2;
  assign mem[2610] = 9'd3;
  assign mem[2611] = 9'd4;
  assign mem[2612] = 9'd5;
  assign mem[2613] = 9'd6;
  assign mem[2614] = 9'd7;
  assign mem[2615] = 9'd8;
  assign mem[2616] = 9'd2;
  assign mem[2617] = 9'd3;
  assign mem[2618] = 9'd4;
  assign mem[2619] = 9'd5;
  assign mem[2620] = 9'd6;
  assign mem[2621] = 9'd7;
  assign mem[2622] = 9'd8;
  assign mem[2623] = 9'd9;
  assign mem[2624] = 9'd6;
  assign mem[2625] = 9'd5;
  assign mem[2626] = 9'd6;
  assign mem[2627] = 9'd7;
  assign mem[2628] = 9'd8;
  assign mem[2629] = 9'd9;
  assign mem[2630] = 9'd10;
  assign mem[2631] = 9'd11;
  assign mem[2632] = 9'd5;
  assign mem[2633] = 9'd4;
  assign mem[2634] = 9'd5;
  assign mem[2635] = 9'd6;
  assign mem[2636] = 9'd7;
  assign mem[2637] = 9'd8;
  assign mem[2638] = 9'd9;
  assign mem[2639] = 9'd10;
  assign mem[2640] = 9'd4;
  assign mem[2641] = 9'd3;
  assign mem[2642] = 9'd4;
  assign mem[2643] = 9'd5;
  assign mem[2644] = 9'd6;
  assign mem[2645] = 9'd7;
  assign mem[2646] = 9'd8;
  assign mem[2647] = 9'd9;
  assign mem[2648] = 9'd3;
  assign mem[2649] = 9'd2;
  assign mem[2650] = 9'd3;
  assign mem[2651] = 9'd4;
  assign mem[2652] = 9'd5;
  assign mem[2653] = 9'd6;
  assign mem[2654] = 9'd7;
  assign mem[2655] = 9'd8;
  assign mem[2656] = 9'd2;
  assign mem[2657] = 9'd1;
  assign mem[2658] = 9'd2;
  assign mem[2659] = 9'd3;
  assign mem[2660] = 9'd4;
  assign mem[2661] = 9'd5;
  assign mem[2662] = 9'd6;
  assign mem[2663] = 9'd7;
  assign mem[2664] = 9'd1;
  assign mem[2665] = 9'd0;
  assign mem[2666] = 9'd1;
  assign mem[2667] = 9'd2;
  assign mem[2668] = 9'd3;
  assign mem[2669] = 9'd4;
  assign mem[2670] = 9'd5;
  assign mem[2671] = 9'd6;
  assign mem[2672] = 9'd2;
  assign mem[2673] = 9'd1;
  assign mem[2674] = 9'd2;
  assign mem[2675] = 9'd3;
  assign mem[2676] = 9'd4;
  assign mem[2677] = 9'd5;
  assign mem[2678] = 9'd6;
  assign mem[2679] = 9'd7;
  assign mem[2680] = 9'd3;
  assign mem[2681] = 9'd2;
  assign mem[2682] = 9'd3;
  assign mem[2683] = 9'd4;
  assign mem[2684] = 9'd5;
  assign mem[2685] = 9'd6;
  assign mem[2686] = 9'd7;
  assign mem[2687] = 9'd8;
  assign mem[2688] = 9'd7;
  assign mem[2689] = 9'd6;
  assign mem[2690] = 9'd5;
  assign mem[2691] = 9'd6;
  assign mem[2692] = 9'd7;
  assign mem[2693] = 9'd8;
  assign mem[2694] = 9'd9;
  assign mem[2695] = 9'd10;
  assign mem[2696] = 9'd6;
  assign mem[2697] = 9'd5;
  assign mem[2698] = 9'd4;
  assign mem[2699] = 9'd5;
  assign mem[2700] = 9'd6;
  assign mem[2701] = 9'd7;
  assign mem[2702] = 9'd8;
  assign mem[2703] = 9'd9;
  assign mem[2704] = 9'd5;
  assign mem[2705] = 9'd4;
  assign mem[2706] = 9'd3;
  assign mem[2707] = 9'd4;
  assign mem[2708] = 9'd5;
  assign mem[2709] = 9'd6;
  assign mem[2710] = 9'd7;
  assign mem[2711] = 9'd8;
  assign mem[2712] = 9'd4;
  assign mem[2713] = 9'd3;
  assign mem[2714] = 9'd2;
  assign mem[2715] = 9'd3;
  assign mem[2716] = 9'd4;
  assign mem[2717] = 9'd5;
  assign mem[2718] = 9'd6;
  assign mem[2719] = 9'd7;
  assign mem[2720] = 9'd3;
  assign mem[2721] = 9'd2;
  assign mem[2722] = 9'd1;
  assign mem[2723] = 9'd2;
  assign mem[2724] = 9'd3;
  assign mem[2725] = 9'd4;
  assign mem[2726] = 9'd5;
  assign mem[2727] = 9'd6;
  assign mem[2728] = 9'd2;
  assign mem[2729] = 9'd1;
  assign mem[2730] = 9'd0;
  assign mem[2731] = 9'd1;
  assign mem[2732] = 9'd2;
  assign mem[2733] = 9'd3;
  assign mem[2734] = 9'd4;
  assign mem[2735] = 9'd5;
  assign mem[2736] = 9'd3;
  assign mem[2737] = 9'd2;
  assign mem[2738] = 9'd1;
  assign mem[2739] = 9'd2;
  assign mem[2740] = 9'd3;
  assign mem[2741] = 9'd4;
  assign mem[2742] = 9'd5;
  assign mem[2743] = 9'd6;
  assign mem[2744] = 9'd4;
  assign mem[2745] = 9'd3;
  assign mem[2746] = 9'd2;
  assign mem[2747] = 9'd3;
  assign mem[2748] = 9'd4;
  assign mem[2749] = 9'd5;
  assign mem[2750] = 9'd6;
  assign mem[2751] = 9'd7;
  assign mem[2752] = 9'd8;
  assign mem[2753] = 9'd7;
  assign mem[2754] = 9'd6;
  assign mem[2755] = 9'd5;
  assign mem[2756] = 9'd6;
  assign mem[2757] = 9'd7;
  assign mem[2758] = 9'd8;
  assign mem[2759] = 9'd9;
  assign mem[2760] = 9'd7;
  assign mem[2761] = 9'd6;
  assign mem[2762] = 9'd5;
  assign mem[2763] = 9'd4;
  assign mem[2764] = 9'd5;
  assign mem[2765] = 9'd6;
  assign mem[2766] = 9'd7;
  assign mem[2767] = 9'd8;
  assign mem[2768] = 9'd6;
  assign mem[2769] = 9'd5;
  assign mem[2770] = 9'd4;
  assign mem[2771] = 9'd3;
  assign mem[2772] = 9'd4;
  assign mem[2773] = 9'd5;
  assign mem[2774] = 9'd6;
  assign mem[2775] = 9'd7;
  assign mem[2776] = 9'd5;
  assign mem[2777] = 9'd4;
  assign mem[2778] = 9'd3;
  assign mem[2779] = 9'd2;
  assign mem[2780] = 9'd3;
  assign mem[2781] = 9'd4;
  assign mem[2782] = 9'd5;
  assign mem[2783] = 9'd6;
  assign mem[2784] = 9'd4;
  assign mem[2785] = 9'd3;
  assign mem[2786] = 9'd2;
  assign mem[2787] = 9'd1;
  assign mem[2788] = 9'd2;
  assign mem[2789] = 9'd3;
  assign mem[2790] = 9'd4;
  assign mem[2791] = 9'd5;
  assign mem[2792] = 9'd3;
  assign mem[2793] = 9'd2;
  assign mem[2794] = 9'd1;
  assign mem[2795] = 9'd0;
  assign mem[2796] = 9'd1;
  assign mem[2797] = 9'd2;
  assign mem[2798] = 9'd3;
  assign mem[2799] = 9'd4;
  assign mem[2800] = 9'd4;
  assign mem[2801] = 9'd3;
  assign mem[2802] = 9'd2;
  assign mem[2803] = 9'd1;
  assign mem[2804] = 9'd2;
  assign mem[2805] = 9'd3;
  assign mem[2806] = 9'd4;
  assign mem[2807] = 9'd5;
  assign mem[2808] = 9'd5;
  assign mem[2809] = 9'd4;
  assign mem[2810] = 9'd3;
  assign mem[2811] = 9'd2;
  assign mem[2812] = 9'd3;
  assign mem[2813] = 9'd4;
  assign mem[2814] = 9'd5;
  assign mem[2815] = 9'd6;
  assign mem[2816] = 9'd9;
  assign mem[2817] = 9'd8;
  assign mem[2818] = 9'd7;
  assign mem[2819] = 9'd6;
  assign mem[2820] = 9'd5;
  assign mem[2821] = 9'd6;
  assign mem[2822] = 9'd7;
  assign mem[2823] = 9'd8;
  assign mem[2824] = 9'd8;
  assign mem[2825] = 9'd7;
  assign mem[2826] = 9'd6;
  assign mem[2827] = 9'd5;
  assign mem[2828] = 9'd4;
  assign mem[2829] = 9'd5;
  assign mem[2830] = 9'd6;
  assign mem[2831] = 9'd7;
  assign mem[2832] = 9'd7;
  assign mem[2833] = 9'd6;
  assign mem[2834] = 9'd5;
  assign mem[2835] = 9'd4;
  assign mem[2836] = 9'd3;
  assign mem[2837] = 9'd4;
  assign mem[2838] = 9'd5;
  assign mem[2839] = 9'd6;
  assign mem[2840] = 9'd6;
  assign mem[2841] = 9'd5;
  assign mem[2842] = 9'd4;
  assign mem[2843] = 9'd3;
  assign mem[2844] = 9'd2;
  assign mem[2845] = 9'd3;
  assign mem[2846] = 9'd4;
  assign mem[2847] = 9'd5;
  assign mem[2848] = 9'd5;
  assign mem[2849] = 9'd4;
  assign mem[2850] = 9'd3;
  assign mem[2851] = 9'd2;
  assign mem[2852] = 9'd1;
  assign mem[2853] = 9'd2;
  assign mem[2854] = 9'd3;
  assign mem[2855] = 9'd4;
  assign mem[2856] = 9'd4;
  assign mem[2857] = 9'd3;
  assign mem[2858] = 9'd2;
  assign mem[2859] = 9'd1;
  assign mem[2860] = 9'd0;
  assign mem[2861] = 9'd1;
  assign mem[2862] = 9'd2;
  assign mem[2863] = 9'd3;
  assign mem[2864] = 9'd5;
  assign mem[2865] = 9'd4;
  assign mem[2866] = 9'd3;
  assign mem[2867] = 9'd2;
  assign mem[2868] = 9'd1;
  assign mem[2869] = 9'd2;
  assign mem[2870] = 9'd3;
  assign mem[2871] = 9'd4;
  assign mem[2872] = 9'd6;
  assign mem[2873] = 9'd5;
  assign mem[2874] = 9'd4;
  assign mem[2875] = 9'd3;
  assign mem[2876] = 9'd2;
  assign mem[2877] = 9'd3;
  assign mem[2878] = 9'd4;
  assign mem[2879] = 9'd5;
  assign mem[2880] = 9'd10;
  assign mem[2881] = 9'd9;
  assign mem[2882] = 9'd8;
  assign mem[2883] = 9'd7;
  assign mem[2884] = 9'd6;
  assign mem[2885] = 9'd5;
  assign mem[2886] = 9'd6;
  assign mem[2887] = 9'd7;
  assign mem[2888] = 9'd9;
  assign mem[2889] = 9'd8;
  assign mem[2890] = 9'd7;
  assign mem[2891] = 9'd6;
  assign mem[2892] = 9'd5;
  assign mem[2893] = 9'd4;
  assign mem[2894] = 9'd5;
  assign mem[2895] = 9'd6;
  assign mem[2896] = 9'd8;
  assign mem[2897] = 9'd7;
  assign mem[2898] = 9'd6;
  assign mem[2899] = 9'd5;
  assign mem[2900] = 9'd4;
  assign mem[2901] = 9'd3;
  assign mem[2902] = 9'd4;
  assign mem[2903] = 9'd5;
  assign mem[2904] = 9'd7;
  assign mem[2905] = 9'd6;
  assign mem[2906] = 9'd5;
  assign mem[2907] = 9'd4;
  assign mem[2908] = 9'd3;
  assign mem[2909] = 9'd2;
  assign mem[2910] = 9'd3;
  assign mem[2911] = 9'd4;
  assign mem[2912] = 9'd6;
  assign mem[2913] = 9'd5;
  assign mem[2914] = 9'd4;
  assign mem[2915] = 9'd3;
  assign mem[2916] = 9'd2;
  assign mem[2917] = 9'd1;
  assign mem[2918] = 9'd2;
  assign mem[2919] = 9'd3;
  assign mem[2920] = 9'd5;
  assign mem[2921] = 9'd4;
  assign mem[2922] = 9'd3;
  assign mem[2923] = 9'd2;
  assign mem[2924] = 9'd1;
  assign mem[2925] = 9'd0;
  assign mem[2926] = 9'd1;
  assign mem[2927] = 9'd2;
  assign mem[2928] = 9'd6;
  assign mem[2929] = 9'd5;
  assign mem[2930] = 9'd4;
  assign mem[2931] = 9'd3;
  assign mem[2932] = 9'd2;
  assign mem[2933] = 9'd1;
  assign mem[2934] = 9'd2;
  assign mem[2935] = 9'd3;
  assign mem[2936] = 9'd7;
  assign mem[2937] = 9'd6;
  assign mem[2938] = 9'd5;
  assign mem[2939] = 9'd4;
  assign mem[2940] = 9'd3;
  assign mem[2941] = 9'd2;
  assign mem[2942] = 9'd3;
  assign mem[2943] = 9'd4;
  assign mem[2944] = 9'd11;
  assign mem[2945] = 9'd10;
  assign mem[2946] = 9'd9;
  assign mem[2947] = 9'd8;
  assign mem[2948] = 9'd7;
  assign mem[2949] = 9'd6;
  assign mem[2950] = 9'd5;
  assign mem[2951] = 9'd6;
  assign mem[2952] = 9'd10;
  assign mem[2953] = 9'd9;
  assign mem[2954] = 9'd8;
  assign mem[2955] = 9'd7;
  assign mem[2956] = 9'd6;
  assign mem[2957] = 9'd5;
  assign mem[2958] = 9'd4;
  assign mem[2959] = 9'd5;
  assign mem[2960] = 9'd9;
  assign mem[2961] = 9'd8;
  assign mem[2962] = 9'd7;
  assign mem[2963] = 9'd6;
  assign mem[2964] = 9'd5;
  assign mem[2965] = 9'd4;
  assign mem[2966] = 9'd3;
  assign mem[2967] = 9'd4;
  assign mem[2968] = 9'd8;
  assign mem[2969] = 9'd7;
  assign mem[2970] = 9'd6;
  assign mem[2971] = 9'd5;
  assign mem[2972] = 9'd4;
  assign mem[2973] = 9'd3;
  assign mem[2974] = 9'd2;
  assign mem[2975] = 9'd3;
  assign mem[2976] = 9'd7;
  assign mem[2977] = 9'd6;
  assign mem[2978] = 9'd5;
  assign mem[2979] = 9'd4;
  assign mem[2980] = 9'd3;
  assign mem[2981] = 9'd2;
  assign mem[2982] = 9'd1;
  assign mem[2983] = 9'd2;
  assign mem[2984] = 9'd6;
  assign mem[2985] = 9'd5;
  assign mem[2986] = 9'd4;
  assign mem[2987] = 9'd3;
  assign mem[2988] = 9'd2;
  assign mem[2989] = 9'd1;
  assign mem[2990] = 9'd0;
  assign mem[2991] = 9'd1;
  assign mem[2992] = 9'd7;
  assign mem[2993] = 9'd6;
  assign mem[2994] = 9'd5;
  assign mem[2995] = 9'd4;
  assign mem[2996] = 9'd3;
  assign mem[2997] = 9'd2;
  assign mem[2998] = 9'd1;
  assign mem[2999] = 9'd2;
  assign mem[3000] = 9'd8;
  assign mem[3001] = 9'd7;
  assign mem[3002] = 9'd6;
  assign mem[3003] = 9'd5;
  assign mem[3004] = 9'd4;
  assign mem[3005] = 9'd3;
  assign mem[3006] = 9'd2;
  assign mem[3007] = 9'd3;
  assign mem[3008] = 9'd12;
  assign mem[3009] = 9'd11;
  assign mem[3010] = 9'd10;
  assign mem[3011] = 9'd9;
  assign mem[3012] = 9'd8;
  assign mem[3013] = 9'd7;
  assign mem[3014] = 9'd6;
  assign mem[3015] = 9'd5;
  assign mem[3016] = 9'd11;
  assign mem[3017] = 9'd10;
  assign mem[3018] = 9'd9;
  assign mem[3019] = 9'd8;
  assign mem[3020] = 9'd7;
  assign mem[3021] = 9'd6;
  assign mem[3022] = 9'd5;
  assign mem[3023] = 9'd4;
  assign mem[3024] = 9'd10;
  assign mem[3025] = 9'd9;
  assign mem[3026] = 9'd8;
  assign mem[3027] = 9'd7;
  assign mem[3028] = 9'd6;
  assign mem[3029] = 9'd5;
  assign mem[3030] = 9'd4;
  assign mem[3031] = 9'd3;
  assign mem[3032] = 9'd9;
  assign mem[3033] = 9'd8;
  assign mem[3034] = 9'd7;
  assign mem[3035] = 9'd6;
  assign mem[3036] = 9'd5;
  assign mem[3037] = 9'd4;
  assign mem[3038] = 9'd3;
  assign mem[3039] = 9'd2;
  assign mem[3040] = 9'd8;
  assign mem[3041] = 9'd7;
  assign mem[3042] = 9'd6;
  assign mem[3043] = 9'd5;
  assign mem[3044] = 9'd4;
  assign mem[3045] = 9'd3;
  assign mem[3046] = 9'd2;
  assign mem[3047] = 9'd1;
  assign mem[3048] = 9'd7;
  assign mem[3049] = 9'd6;
  assign mem[3050] = 9'd5;
  assign mem[3051] = 9'd4;
  assign mem[3052] = 9'd3;
  assign mem[3053] = 9'd2;
  assign mem[3054] = 9'd1;
  assign mem[3055] = 9'd0;
  assign mem[3056] = 9'd8;
  assign mem[3057] = 9'd7;
  assign mem[3058] = 9'd6;
  assign mem[3059] = 9'd5;
  assign mem[3060] = 9'd4;
  assign mem[3061] = 9'd3;
  assign mem[3062] = 9'd2;
  assign mem[3063] = 9'd1;
  assign mem[3064] = 9'd9;
  assign mem[3065] = 9'd8;
  assign mem[3066] = 9'd7;
  assign mem[3067] = 9'd6;
  assign mem[3068] = 9'd5;
  assign mem[3069] = 9'd4;
  assign mem[3070] = 9'd3;
  assign mem[3071] = 9'd2;
  assign mem[3072] = 9'd6;
  assign mem[3073] = 9'd7;
  assign mem[3074] = 9'd8;
  assign mem[3075] = 9'd9;
  assign mem[3076] = 9'd10;
  assign mem[3077] = 9'd11;
  assign mem[3078] = 9'd12;
  assign mem[3079] = 9'd13;
  assign mem[3080] = 9'd5;
  assign mem[3081] = 9'd6;
  assign mem[3082] = 9'd7;
  assign mem[3083] = 9'd8;
  assign mem[3084] = 9'd9;
  assign mem[3085] = 9'd10;
  assign mem[3086] = 9'd11;
  assign mem[3087] = 9'd12;
  assign mem[3088] = 9'd4;
  assign mem[3089] = 9'd5;
  assign mem[3090] = 9'd6;
  assign mem[3091] = 9'd7;
  assign mem[3092] = 9'd8;
  assign mem[3093] = 9'd9;
  assign mem[3094] = 9'd10;
  assign mem[3095] = 9'd11;
  assign mem[3096] = 9'd3;
  assign mem[3097] = 9'd4;
  assign mem[3098] = 9'd5;
  assign mem[3099] = 9'd6;
  assign mem[3100] = 9'd7;
  assign mem[3101] = 9'd8;
  assign mem[3102] = 9'd9;
  assign mem[3103] = 9'd10;
  assign mem[3104] = 9'd2;
  assign mem[3105] = 9'd3;
  assign mem[3106] = 9'd4;
  assign mem[3107] = 9'd5;
  assign mem[3108] = 9'd6;
  assign mem[3109] = 9'd7;
  assign mem[3110] = 9'd8;
  assign mem[3111] = 9'd9;
  assign mem[3112] = 9'd1;
  assign mem[3113] = 9'd2;
  assign mem[3114] = 9'd3;
  assign mem[3115] = 9'd4;
  assign mem[3116] = 9'd5;
  assign mem[3117] = 9'd6;
  assign mem[3118] = 9'd7;
  assign mem[3119] = 9'd8;
  assign mem[3120] = 9'd0;
  assign mem[3121] = 9'd1;
  assign mem[3122] = 9'd2;
  assign mem[3123] = 9'd3;
  assign mem[3124] = 9'd4;
  assign mem[3125] = 9'd5;
  assign mem[3126] = 9'd6;
  assign mem[3127] = 9'd7;
  assign mem[3128] = 9'd1;
  assign mem[3129] = 9'd2;
  assign mem[3130] = 9'd3;
  assign mem[3131] = 9'd4;
  assign mem[3132] = 9'd5;
  assign mem[3133] = 9'd6;
  assign mem[3134] = 9'd7;
  assign mem[3135] = 9'd8;
  assign mem[3136] = 9'd7;
  assign mem[3137] = 9'd6;
  assign mem[3138] = 9'd7;
  assign mem[3139] = 9'd8;
  assign mem[3140] = 9'd9;
  assign mem[3141] = 9'd10;
  assign mem[3142] = 9'd11;
  assign mem[3143] = 9'd12;
  assign mem[3144] = 9'd6;
  assign mem[3145] = 9'd5;
  assign mem[3146] = 9'd6;
  assign mem[3147] = 9'd7;
  assign mem[3148] = 9'd8;
  assign mem[3149] = 9'd9;
  assign mem[3150] = 9'd10;
  assign mem[3151] = 9'd11;
  assign mem[3152] = 9'd5;
  assign mem[3153] = 9'd4;
  assign mem[3154] = 9'd5;
  assign mem[3155] = 9'd6;
  assign mem[3156] = 9'd7;
  assign mem[3157] = 9'd8;
  assign mem[3158] = 9'd9;
  assign mem[3159] = 9'd10;
  assign mem[3160] = 9'd4;
  assign mem[3161] = 9'd3;
  assign mem[3162] = 9'd4;
  assign mem[3163] = 9'd5;
  assign mem[3164] = 9'd6;
  assign mem[3165] = 9'd7;
  assign mem[3166] = 9'd8;
  assign mem[3167] = 9'd9;
  assign mem[3168] = 9'd3;
  assign mem[3169] = 9'd2;
  assign mem[3170] = 9'd3;
  assign mem[3171] = 9'd4;
  assign mem[3172] = 9'd5;
  assign mem[3173] = 9'd6;
  assign mem[3174] = 9'd7;
  assign mem[3175] = 9'd8;
  assign mem[3176] = 9'd2;
  assign mem[3177] = 9'd1;
  assign mem[3178] = 9'd2;
  assign mem[3179] = 9'd3;
  assign mem[3180] = 9'd4;
  assign mem[3181] = 9'd5;
  assign mem[3182] = 9'd6;
  assign mem[3183] = 9'd7;
  assign mem[3184] = 9'd1;
  assign mem[3185] = 9'd0;
  assign mem[3186] = 9'd1;
  assign mem[3187] = 9'd2;
  assign mem[3188] = 9'd3;
  assign mem[3189] = 9'd4;
  assign mem[3190] = 9'd5;
  assign mem[3191] = 9'd6;
  assign mem[3192] = 9'd2;
  assign mem[3193] = 9'd1;
  assign mem[3194] = 9'd2;
  assign mem[3195] = 9'd3;
  assign mem[3196] = 9'd4;
  assign mem[3197] = 9'd5;
  assign mem[3198] = 9'd6;
  assign mem[3199] = 9'd7;
  assign mem[3200] = 9'd8;
  assign mem[3201] = 9'd7;
  assign mem[3202] = 9'd6;
  assign mem[3203] = 9'd7;
  assign mem[3204] = 9'd8;
  assign mem[3205] = 9'd9;
  assign mem[3206] = 9'd10;
  assign mem[3207] = 9'd11;
  assign mem[3208] = 9'd7;
  assign mem[3209] = 9'd6;
  assign mem[3210] = 9'd5;
  assign mem[3211] = 9'd6;
  assign mem[3212] = 9'd7;
  assign mem[3213] = 9'd8;
  assign mem[3214] = 9'd9;
  assign mem[3215] = 9'd10;
  assign mem[3216] = 9'd6;
  assign mem[3217] = 9'd5;
  assign mem[3218] = 9'd4;
  assign mem[3219] = 9'd5;
  assign mem[3220] = 9'd6;
  assign mem[3221] = 9'd7;
  assign mem[3222] = 9'd8;
  assign mem[3223] = 9'd9;
  assign mem[3224] = 9'd5;
  assign mem[3225] = 9'd4;
  assign mem[3226] = 9'd3;
  assign mem[3227] = 9'd4;
  assign mem[3228] = 9'd5;
  assign mem[3229] = 9'd6;
  assign mem[3230] = 9'd7;
  assign mem[3231] = 9'd8;
  assign mem[3232] = 9'd4;
  assign mem[3233] = 9'd3;
  assign mem[3234] = 9'd2;
  assign mem[3235] = 9'd3;
  assign mem[3236] = 9'd4;
  assign mem[3237] = 9'd5;
  assign mem[3238] = 9'd6;
  assign mem[3239] = 9'd7;
  assign mem[3240] = 9'd3;
  assign mem[3241] = 9'd2;
  assign mem[3242] = 9'd1;
  assign mem[3243] = 9'd2;
  assign mem[3244] = 9'd3;
  assign mem[3245] = 9'd4;
  assign mem[3246] = 9'd5;
  assign mem[3247] = 9'd6;
  assign mem[3248] = 9'd2;
  assign mem[3249] = 9'd1;
  assign mem[3250] = 9'd0;
  assign mem[3251] = 9'd1;
  assign mem[3252] = 9'd2;
  assign mem[3253] = 9'd3;
  assign mem[3254] = 9'd4;
  assign mem[3255] = 9'd5;
  assign mem[3256] = 9'd3;
  assign mem[3257] = 9'd2;
  assign mem[3258] = 9'd1;
  assign mem[3259] = 9'd2;
  assign mem[3260] = 9'd3;
  assign mem[3261] = 9'd4;
  assign mem[3262] = 9'd5;
  assign mem[3263] = 9'd6;
  assign mem[3264] = 9'd9;
  assign mem[3265] = 9'd8;
  assign mem[3266] = 9'd7;
  assign mem[3267] = 9'd6;
  assign mem[3268] = 9'd7;
  assign mem[3269] = 9'd8;
  assign mem[3270] = 9'd9;
  assign mem[3271] = 9'd10;
  assign mem[3272] = 9'd8;
  assign mem[3273] = 9'd7;
  assign mem[3274] = 9'd6;
  assign mem[3275] = 9'd5;
  assign mem[3276] = 9'd6;
  assign mem[3277] = 9'd7;
  assign mem[3278] = 9'd8;
  assign mem[3279] = 9'd9;
  assign mem[3280] = 9'd7;
  assign mem[3281] = 9'd6;
  assign mem[3282] = 9'd5;
  assign mem[3283] = 9'd4;
  assign mem[3284] = 9'd5;
  assign mem[3285] = 9'd6;
  assign mem[3286] = 9'd7;
  assign mem[3287] = 9'd8;
  assign mem[3288] = 9'd6;
  assign mem[3289] = 9'd5;
  assign mem[3290] = 9'd4;
  assign mem[3291] = 9'd3;
  assign mem[3292] = 9'd4;
  assign mem[3293] = 9'd5;
  assign mem[3294] = 9'd6;
  assign mem[3295] = 9'd7;
  assign mem[3296] = 9'd5;
  assign mem[3297] = 9'd4;
  assign mem[3298] = 9'd3;
  assign mem[3299] = 9'd2;
  assign mem[3300] = 9'd3;
  assign mem[3301] = 9'd4;
  assign mem[3302] = 9'd5;
  assign mem[3303] = 9'd6;
  assign mem[3304] = 9'd4;
  assign mem[3305] = 9'd3;
  assign mem[3306] = 9'd2;
  assign mem[3307] = 9'd1;
  assign mem[3308] = 9'd2;
  assign mem[3309] = 9'd3;
  assign mem[3310] = 9'd4;
  assign mem[3311] = 9'd5;
  assign mem[3312] = 9'd3;
  assign mem[3313] = 9'd2;
  assign mem[3314] = 9'd1;
  assign mem[3315] = 9'd0;
  assign mem[3316] = 9'd1;
  assign mem[3317] = 9'd2;
  assign mem[3318] = 9'd3;
  assign mem[3319] = 9'd4;
  assign mem[3320] = 9'd4;
  assign mem[3321] = 9'd3;
  assign mem[3322] = 9'd2;
  assign mem[3323] = 9'd1;
  assign mem[3324] = 9'd2;
  assign mem[3325] = 9'd3;
  assign mem[3326] = 9'd4;
  assign mem[3327] = 9'd5;
  assign mem[3328] = 9'd10;
  assign mem[3329] = 9'd9;
  assign mem[3330] = 9'd8;
  assign mem[3331] = 9'd7;
  assign mem[3332] = 9'd6;
  assign mem[3333] = 9'd7;
  assign mem[3334] = 9'd8;
  assign mem[3335] = 9'd9;
  assign mem[3336] = 9'd9;
  assign mem[3337] = 9'd8;
  assign mem[3338] = 9'd7;
  assign mem[3339] = 9'd6;
  assign mem[3340] = 9'd5;
  assign mem[3341] = 9'd6;
  assign mem[3342] = 9'd7;
  assign mem[3343] = 9'd8;
  assign mem[3344] = 9'd8;
  assign mem[3345] = 9'd7;
  assign mem[3346] = 9'd6;
  assign mem[3347] = 9'd5;
  assign mem[3348] = 9'd4;
  assign mem[3349] = 9'd5;
  assign mem[3350] = 9'd6;
  assign mem[3351] = 9'd7;
  assign mem[3352] = 9'd7;
  assign mem[3353] = 9'd6;
  assign mem[3354] = 9'd5;
  assign mem[3355] = 9'd4;
  assign mem[3356] = 9'd3;
  assign mem[3357] = 9'd4;
  assign mem[3358] = 9'd5;
  assign mem[3359] = 9'd6;
  assign mem[3360] = 9'd6;
  assign mem[3361] = 9'd5;
  assign mem[3362] = 9'd4;
  assign mem[3363] = 9'd3;
  assign mem[3364] = 9'd2;
  assign mem[3365] = 9'd3;
  assign mem[3366] = 9'd4;
  assign mem[3367] = 9'd5;
  assign mem[3368] = 9'd5;
  assign mem[3369] = 9'd4;
  assign mem[3370] = 9'd3;
  assign mem[3371] = 9'd2;
  assign mem[3372] = 9'd1;
  assign mem[3373] = 9'd2;
  assign mem[3374] = 9'd3;
  assign mem[3375] = 9'd4;
  assign mem[3376] = 9'd4;
  assign mem[3377] = 9'd3;
  assign mem[3378] = 9'd2;
  assign mem[3379] = 9'd1;
  assign mem[3380] = 9'd0;
  assign mem[3381] = 9'd1;
  assign mem[3382] = 9'd2;
  assign mem[3383] = 9'd3;
  assign mem[3384] = 9'd5;
  assign mem[3385] = 9'd4;
  assign mem[3386] = 9'd3;
  assign mem[3387] = 9'd2;
  assign mem[3388] = 9'd1;
  assign mem[3389] = 9'd2;
  assign mem[3390] = 9'd3;
  assign mem[3391] = 9'd4;
  assign mem[3392] = 9'd11;
  assign mem[3393] = 9'd10;
  assign mem[3394] = 9'd9;
  assign mem[3395] = 9'd8;
  assign mem[3396] = 9'd7;
  assign mem[3397] = 9'd6;
  assign mem[3398] = 9'd7;
  assign mem[3399] = 9'd8;
  assign mem[3400] = 9'd10;
  assign mem[3401] = 9'd9;
  assign mem[3402] = 9'd8;
  assign mem[3403] = 9'd7;
  assign mem[3404] = 9'd6;
  assign mem[3405] = 9'd5;
  assign mem[3406] = 9'd6;
  assign mem[3407] = 9'd7;
  assign mem[3408] = 9'd9;
  assign mem[3409] = 9'd8;
  assign mem[3410] = 9'd7;
  assign mem[3411] = 9'd6;
  assign mem[3412] = 9'd5;
  assign mem[3413] = 9'd4;
  assign mem[3414] = 9'd5;
  assign mem[3415] = 9'd6;
  assign mem[3416] = 9'd8;
  assign mem[3417] = 9'd7;
  assign mem[3418] = 9'd6;
  assign mem[3419] = 9'd5;
  assign mem[3420] = 9'd4;
  assign mem[3421] = 9'd3;
  assign mem[3422] = 9'd4;
  assign mem[3423] = 9'd5;
  assign mem[3424] = 9'd7;
  assign mem[3425] = 9'd6;
  assign mem[3426] = 9'd5;
  assign mem[3427] = 9'd4;
  assign mem[3428] = 9'd3;
  assign mem[3429] = 9'd2;
  assign mem[3430] = 9'd3;
  assign mem[3431] = 9'd4;
  assign mem[3432] = 9'd6;
  assign mem[3433] = 9'd5;
  assign mem[3434] = 9'd4;
  assign mem[3435] = 9'd3;
  assign mem[3436] = 9'd2;
  assign mem[3437] = 9'd1;
  assign mem[3438] = 9'd2;
  assign mem[3439] = 9'd3;
  assign mem[3440] = 9'd5;
  assign mem[3441] = 9'd4;
  assign mem[3442] = 9'd3;
  assign mem[3443] = 9'd2;
  assign mem[3444] = 9'd1;
  assign mem[3445] = 9'd0;
  assign mem[3446] = 9'd1;
  assign mem[3447] = 9'd2;
  assign mem[3448] = 9'd6;
  assign mem[3449] = 9'd5;
  assign mem[3450] = 9'd4;
  assign mem[3451] = 9'd3;
  assign mem[3452] = 9'd2;
  assign mem[3453] = 9'd1;
  assign mem[3454] = 9'd2;
  assign mem[3455] = 9'd3;
  assign mem[3456] = 9'd12;
  assign mem[3457] = 9'd11;
  assign mem[3458] = 9'd10;
  assign mem[3459] = 9'd9;
  assign mem[3460] = 9'd8;
  assign mem[3461] = 9'd7;
  assign mem[3462] = 9'd6;
  assign mem[3463] = 9'd7;
  assign mem[3464] = 9'd11;
  assign mem[3465] = 9'd10;
  assign mem[3466] = 9'd9;
  assign mem[3467] = 9'd8;
  assign mem[3468] = 9'd7;
  assign mem[3469] = 9'd6;
  assign mem[3470] = 9'd5;
  assign mem[3471] = 9'd6;
  assign mem[3472] = 9'd10;
  assign mem[3473] = 9'd9;
  assign mem[3474] = 9'd8;
  assign mem[3475] = 9'd7;
  assign mem[3476] = 9'd6;
  assign mem[3477] = 9'd5;
  assign mem[3478] = 9'd4;
  assign mem[3479] = 9'd5;
  assign mem[3480] = 9'd9;
  assign mem[3481] = 9'd8;
  assign mem[3482] = 9'd7;
  assign mem[3483] = 9'd6;
  assign mem[3484] = 9'd5;
  assign mem[3485] = 9'd4;
  assign mem[3486] = 9'd3;
  assign mem[3487] = 9'd4;
  assign mem[3488] = 9'd8;
  assign mem[3489] = 9'd7;
  assign mem[3490] = 9'd6;
  assign mem[3491] = 9'd5;
  assign mem[3492] = 9'd4;
  assign mem[3493] = 9'd3;
  assign mem[3494] = 9'd2;
  assign mem[3495] = 9'd3;
  assign mem[3496] = 9'd7;
  assign mem[3497] = 9'd6;
  assign mem[3498] = 9'd5;
  assign mem[3499] = 9'd4;
  assign mem[3500] = 9'd3;
  assign mem[3501] = 9'd2;
  assign mem[3502] = 9'd1;
  assign mem[3503] = 9'd2;
  assign mem[3504] = 9'd6;
  assign mem[3505] = 9'd5;
  assign mem[3506] = 9'd4;
  assign mem[3507] = 9'd3;
  assign mem[3508] = 9'd2;
  assign mem[3509] = 9'd1;
  assign mem[3510] = 9'd0;
  assign mem[3511] = 9'd1;
  assign mem[3512] = 9'd7;
  assign mem[3513] = 9'd6;
  assign mem[3514] = 9'd5;
  assign mem[3515] = 9'd4;
  assign mem[3516] = 9'd3;
  assign mem[3517] = 9'd2;
  assign mem[3518] = 9'd1;
  assign mem[3519] = 9'd2;
  assign mem[3520] = 9'd13;
  assign mem[3521] = 9'd12;
  assign mem[3522] = 9'd11;
  assign mem[3523] = 9'd10;
  assign mem[3524] = 9'd9;
  assign mem[3525] = 9'd8;
  assign mem[3526] = 9'd7;
  assign mem[3527] = 9'd6;
  assign mem[3528] = 9'd12;
  assign mem[3529] = 9'd11;
  assign mem[3530] = 9'd10;
  assign mem[3531] = 9'd9;
  assign mem[3532] = 9'd8;
  assign mem[3533] = 9'd7;
  assign mem[3534] = 9'd6;
  assign mem[3535] = 9'd5;
  assign mem[3536] = 9'd11;
  assign mem[3537] = 9'd10;
  assign mem[3538] = 9'd9;
  assign mem[3539] = 9'd8;
  assign mem[3540] = 9'd7;
  assign mem[3541] = 9'd6;
  assign mem[3542] = 9'd5;
  assign mem[3543] = 9'd4;
  assign mem[3544] = 9'd10;
  assign mem[3545] = 9'd9;
  assign mem[3546] = 9'd8;
  assign mem[3547] = 9'd7;
  assign mem[3548] = 9'd6;
  assign mem[3549] = 9'd5;
  assign mem[3550] = 9'd4;
  assign mem[3551] = 9'd3;
  assign mem[3552] = 9'd9;
  assign mem[3553] = 9'd8;
  assign mem[3554] = 9'd7;
  assign mem[3555] = 9'd6;
  assign mem[3556] = 9'd5;
  assign mem[3557] = 9'd4;
  assign mem[3558] = 9'd3;
  assign mem[3559] = 9'd2;
  assign mem[3560] = 9'd8;
  assign mem[3561] = 9'd7;
  assign mem[3562] = 9'd6;
  assign mem[3563] = 9'd5;
  assign mem[3564] = 9'd4;
  assign mem[3565] = 9'd3;
  assign mem[3566] = 9'd2;
  assign mem[3567] = 9'd1;
  assign mem[3568] = 9'd7;
  assign mem[3569] = 9'd6;
  assign mem[3570] = 9'd5;
  assign mem[3571] = 9'd4;
  assign mem[3572] = 9'd3;
  assign mem[3573] = 9'd2;
  assign mem[3574] = 9'd1;
  assign mem[3575] = 9'd0;
  assign mem[3576] = 9'd8;
  assign mem[3577] = 9'd7;
  assign mem[3578] = 9'd6;
  assign mem[3579] = 9'd5;
  assign mem[3580] = 9'd4;
  assign mem[3581] = 9'd3;
  assign mem[3582] = 9'd2;
  assign mem[3583] = 9'd1;
  assign mem[3584] = 9'd7;
  assign mem[3585] = 9'd8;
  assign mem[3586] = 9'd9;
  assign mem[3587] = 9'd10;
  assign mem[3588] = 9'd11;
  assign mem[3589] = 9'd12;
  assign mem[3590] = 9'd13;
  assign mem[3591] = 9'd14;
  assign mem[3592] = 9'd6;
  assign mem[3593] = 9'd7;
  assign mem[3594] = 9'd8;
  assign mem[3595] = 9'd9;
  assign mem[3596] = 9'd10;
  assign mem[3597] = 9'd11;
  assign mem[3598] = 9'd12;
  assign mem[3599] = 9'd13;
  assign mem[3600] = 9'd5;
  assign mem[3601] = 9'd6;
  assign mem[3602] = 9'd7;
  assign mem[3603] = 9'd8;
  assign mem[3604] = 9'd9;
  assign mem[3605] = 9'd10;
  assign mem[3606] = 9'd11;
  assign mem[3607] = 9'd12;
  assign mem[3608] = 9'd4;
  assign mem[3609] = 9'd5;
  assign mem[3610] = 9'd6;
  assign mem[3611] = 9'd7;
  assign mem[3612] = 9'd8;
  assign mem[3613] = 9'd9;
  assign mem[3614] = 9'd10;
  assign mem[3615] = 9'd11;
  assign mem[3616] = 9'd3;
  assign mem[3617] = 9'd4;
  assign mem[3618] = 9'd5;
  assign mem[3619] = 9'd6;
  assign mem[3620] = 9'd7;
  assign mem[3621] = 9'd8;
  assign mem[3622] = 9'd9;
  assign mem[3623] = 9'd10;
  assign mem[3624] = 9'd2;
  assign mem[3625] = 9'd3;
  assign mem[3626] = 9'd4;
  assign mem[3627] = 9'd5;
  assign mem[3628] = 9'd6;
  assign mem[3629] = 9'd7;
  assign mem[3630] = 9'd8;
  assign mem[3631] = 9'd9;
  assign mem[3632] = 9'd1;
  assign mem[3633] = 9'd2;
  assign mem[3634] = 9'd3;
  assign mem[3635] = 9'd4;
  assign mem[3636] = 9'd5;
  assign mem[3637] = 9'd6;
  assign mem[3638] = 9'd7;
  assign mem[3639] = 9'd8;
  assign mem[3640] = 9'd0;
  assign mem[3641] = 9'd1;
  assign mem[3642] = 9'd2;
  assign mem[3643] = 9'd3;
  assign mem[3644] = 9'd4;
  assign mem[3645] = 9'd5;
  assign mem[3646] = 9'd6;
  assign mem[3647] = 9'd7;
  assign mem[3648] = 9'd8;
  assign mem[3649] = 9'd7;
  assign mem[3650] = 9'd8;
  assign mem[3651] = 9'd9;
  assign mem[3652] = 9'd10;
  assign mem[3653] = 9'd11;
  assign mem[3654] = 9'd12;
  assign mem[3655] = 9'd13;
  assign mem[3656] = 9'd7;
  assign mem[3657] = 9'd6;
  assign mem[3658] = 9'd7;
  assign mem[3659] = 9'd8;
  assign mem[3660] = 9'd9;
  assign mem[3661] = 9'd10;
  assign mem[3662] = 9'd11;
  assign mem[3663] = 9'd12;
  assign mem[3664] = 9'd6;
  assign mem[3665] = 9'd5;
  assign mem[3666] = 9'd6;
  assign mem[3667] = 9'd7;
  assign mem[3668] = 9'd8;
  assign mem[3669] = 9'd9;
  assign mem[3670] = 9'd10;
  assign mem[3671] = 9'd11;
  assign mem[3672] = 9'd5;
  assign mem[3673] = 9'd4;
  assign mem[3674] = 9'd5;
  assign mem[3675] = 9'd6;
  assign mem[3676] = 9'd7;
  assign mem[3677] = 9'd8;
  assign mem[3678] = 9'd9;
  assign mem[3679] = 9'd10;
  assign mem[3680] = 9'd4;
  assign mem[3681] = 9'd3;
  assign mem[3682] = 9'd4;
  assign mem[3683] = 9'd5;
  assign mem[3684] = 9'd6;
  assign mem[3685] = 9'd7;
  assign mem[3686] = 9'd8;
  assign mem[3687] = 9'd9;
  assign mem[3688] = 9'd3;
  assign mem[3689] = 9'd2;
  assign mem[3690] = 9'd3;
  assign mem[3691] = 9'd4;
  assign mem[3692] = 9'd5;
  assign mem[3693] = 9'd6;
  assign mem[3694] = 9'd7;
  assign mem[3695] = 9'd8;
  assign mem[3696] = 9'd2;
  assign mem[3697] = 9'd1;
  assign mem[3698] = 9'd2;
  assign mem[3699] = 9'd3;
  assign mem[3700] = 9'd4;
  assign mem[3701] = 9'd5;
  assign mem[3702] = 9'd6;
  assign mem[3703] = 9'd7;
  assign mem[3704] = 9'd1;
  assign mem[3705] = 9'd0;
  assign mem[3706] = 9'd1;
  assign mem[3707] = 9'd2;
  assign mem[3708] = 9'd3;
  assign mem[3709] = 9'd4;
  assign mem[3710] = 9'd5;
  assign mem[3711] = 9'd6;
  assign mem[3712] = 9'd9;
  assign mem[3713] = 9'd8;
  assign mem[3714] = 9'd7;
  assign mem[3715] = 9'd8;
  assign mem[3716] = 9'd9;
  assign mem[3717] = 9'd10;
  assign mem[3718] = 9'd11;
  assign mem[3719] = 9'd12;
  assign mem[3720] = 9'd8;
  assign mem[3721] = 9'd7;
  assign mem[3722] = 9'd6;
  assign mem[3723] = 9'd7;
  assign mem[3724] = 9'd8;
  assign mem[3725] = 9'd9;
  assign mem[3726] = 9'd10;
  assign mem[3727] = 9'd11;
  assign mem[3728] = 9'd7;
  assign mem[3729] = 9'd6;
  assign mem[3730] = 9'd5;
  assign mem[3731] = 9'd6;
  assign mem[3732] = 9'd7;
  assign mem[3733] = 9'd8;
  assign mem[3734] = 9'd9;
  assign mem[3735] = 9'd10;
  assign mem[3736] = 9'd6;
  assign mem[3737] = 9'd5;
  assign mem[3738] = 9'd4;
  assign mem[3739] = 9'd5;
  assign mem[3740] = 9'd6;
  assign mem[3741] = 9'd7;
  assign mem[3742] = 9'd8;
  assign mem[3743] = 9'd9;
  assign mem[3744] = 9'd5;
  assign mem[3745] = 9'd4;
  assign mem[3746] = 9'd3;
  assign mem[3747] = 9'd4;
  assign mem[3748] = 9'd5;
  assign mem[3749] = 9'd6;
  assign mem[3750] = 9'd7;
  assign mem[3751] = 9'd8;
  assign mem[3752] = 9'd4;
  assign mem[3753] = 9'd3;
  assign mem[3754] = 9'd2;
  assign mem[3755] = 9'd3;
  assign mem[3756] = 9'd4;
  assign mem[3757] = 9'd5;
  assign mem[3758] = 9'd6;
  assign mem[3759] = 9'd7;
  assign mem[3760] = 9'd3;
  assign mem[3761] = 9'd2;
  assign mem[3762] = 9'd1;
  assign mem[3763] = 9'd2;
  assign mem[3764] = 9'd3;
  assign mem[3765] = 9'd4;
  assign mem[3766] = 9'd5;
  assign mem[3767] = 9'd6;
  assign mem[3768] = 9'd2;
  assign mem[3769] = 9'd1;
  assign mem[3770] = 9'd0;
  assign mem[3771] = 9'd1;
  assign mem[3772] = 9'd2;
  assign mem[3773] = 9'd3;
  assign mem[3774] = 9'd4;
  assign mem[3775] = 9'd5;
  assign mem[3776] = 9'd10;
  assign mem[3777] = 9'd9;
  assign mem[3778] = 9'd8;
  assign mem[3779] = 9'd7;
  assign mem[3780] = 9'd8;
  assign mem[3781] = 9'd9;
  assign mem[3782] = 9'd10;
  assign mem[3783] = 9'd11;
  assign mem[3784] = 9'd9;
  assign mem[3785] = 9'd8;
  assign mem[3786] = 9'd7;
  assign mem[3787] = 9'd6;
  assign mem[3788] = 9'd7;
  assign mem[3789] = 9'd8;
  assign mem[3790] = 9'd9;
  assign mem[3791] = 9'd10;
  assign mem[3792] = 9'd8;
  assign mem[3793] = 9'd7;
  assign mem[3794] = 9'd6;
  assign mem[3795] = 9'd5;
  assign mem[3796] = 9'd6;
  assign mem[3797] = 9'd7;
  assign mem[3798] = 9'd8;
  assign mem[3799] = 9'd9;
  assign mem[3800] = 9'd7;
  assign mem[3801] = 9'd6;
  assign mem[3802] = 9'd5;
  assign mem[3803] = 9'd4;
  assign mem[3804] = 9'd5;
  assign mem[3805] = 9'd6;
  assign mem[3806] = 9'd7;
  assign mem[3807] = 9'd8;
  assign mem[3808] = 9'd6;
  assign mem[3809] = 9'd5;
  assign mem[3810] = 9'd4;
  assign mem[3811] = 9'd3;
  assign mem[3812] = 9'd4;
  assign mem[3813] = 9'd5;
  assign mem[3814] = 9'd6;
  assign mem[3815] = 9'd7;
  assign mem[3816] = 9'd5;
  assign mem[3817] = 9'd4;
  assign mem[3818] = 9'd3;
  assign mem[3819] = 9'd2;
  assign mem[3820] = 9'd3;
  assign mem[3821] = 9'd4;
  assign mem[3822] = 9'd5;
  assign mem[3823] = 9'd6;
  assign mem[3824] = 9'd4;
  assign mem[3825] = 9'd3;
  assign mem[3826] = 9'd2;
  assign mem[3827] = 9'd1;
  assign mem[3828] = 9'd2;
  assign mem[3829] = 9'd3;
  assign mem[3830] = 9'd4;
  assign mem[3831] = 9'd5;
  assign mem[3832] = 9'd3;
  assign mem[3833] = 9'd2;
  assign mem[3834] = 9'd1;
  assign mem[3835] = 9'd0;
  assign mem[3836] = 9'd1;
  assign mem[3837] = 9'd2;
  assign mem[3838] = 9'd3;
  assign mem[3839] = 9'd4;
  assign mem[3840] = 9'd11;
  assign mem[3841] = 9'd10;
  assign mem[3842] = 9'd9;
  assign mem[3843] = 9'd8;
  assign mem[3844] = 9'd7;
  assign mem[3845] = 9'd8;
  assign mem[3846] = 9'd9;
  assign mem[3847] = 9'd10;
  assign mem[3848] = 9'd10;
  assign mem[3849] = 9'd9;
  assign mem[3850] = 9'd8;
  assign mem[3851] = 9'd7;
  assign mem[3852] = 9'd6;
  assign mem[3853] = 9'd7;
  assign mem[3854] = 9'd8;
  assign mem[3855] = 9'd9;
  assign mem[3856] = 9'd9;
  assign mem[3857] = 9'd8;
  assign mem[3858] = 9'd7;
  assign mem[3859] = 9'd6;
  assign mem[3860] = 9'd5;
  assign mem[3861] = 9'd6;
  assign mem[3862] = 9'd7;
  assign mem[3863] = 9'd8;
  assign mem[3864] = 9'd8;
  assign mem[3865] = 9'd7;
  assign mem[3866] = 9'd6;
  assign mem[3867] = 9'd5;
  assign mem[3868] = 9'd4;
  assign mem[3869] = 9'd5;
  assign mem[3870] = 9'd6;
  assign mem[3871] = 9'd7;
  assign mem[3872] = 9'd7;
  assign mem[3873] = 9'd6;
  assign mem[3874] = 9'd5;
  assign mem[3875] = 9'd4;
  assign mem[3876] = 9'd3;
  assign mem[3877] = 9'd4;
  assign mem[3878] = 9'd5;
  assign mem[3879] = 9'd6;
  assign mem[3880] = 9'd6;
  assign mem[3881] = 9'd5;
  assign mem[3882] = 9'd4;
  assign mem[3883] = 9'd3;
  assign mem[3884] = 9'd2;
  assign mem[3885] = 9'd3;
  assign mem[3886] = 9'd4;
  assign mem[3887] = 9'd5;
  assign mem[3888] = 9'd5;
  assign mem[3889] = 9'd4;
  assign mem[3890] = 9'd3;
  assign mem[3891] = 9'd2;
  assign mem[3892] = 9'd1;
  assign mem[3893] = 9'd2;
  assign mem[3894] = 9'd3;
  assign mem[3895] = 9'd4;
  assign mem[3896] = 9'd4;
  assign mem[3897] = 9'd3;
  assign mem[3898] = 9'd2;
  assign mem[3899] = 9'd1;
  assign mem[3900] = 9'd0;
  assign mem[3901] = 9'd1;
  assign mem[3902] = 9'd2;
  assign mem[3903] = 9'd3;
  assign mem[3904] = 9'd12;
  assign mem[3905] = 9'd11;
  assign mem[3906] = 9'd10;
  assign mem[3907] = 9'd9;
  assign mem[3908] = 9'd8;
  assign mem[3909] = 9'd7;
  assign mem[3910] = 9'd8;
  assign mem[3911] = 9'd9;
  assign mem[3912] = 9'd11;
  assign mem[3913] = 9'd10;
  assign mem[3914] = 9'd9;
  assign mem[3915] = 9'd8;
  assign mem[3916] = 9'd7;
  assign mem[3917] = 9'd6;
  assign mem[3918] = 9'd7;
  assign mem[3919] = 9'd8;
  assign mem[3920] = 9'd10;
  assign mem[3921] = 9'd9;
  assign mem[3922] = 9'd8;
  assign mem[3923] = 9'd7;
  assign mem[3924] = 9'd6;
  assign mem[3925] = 9'd5;
  assign mem[3926] = 9'd6;
  assign mem[3927] = 9'd7;
  assign mem[3928] = 9'd9;
  assign mem[3929] = 9'd8;
  assign mem[3930] = 9'd7;
  assign mem[3931] = 9'd6;
  assign mem[3932] = 9'd5;
  assign mem[3933] = 9'd4;
  assign mem[3934] = 9'd5;
  assign mem[3935] = 9'd6;
  assign mem[3936] = 9'd8;
  assign mem[3937] = 9'd7;
  assign mem[3938] = 9'd6;
  assign mem[3939] = 9'd5;
  assign mem[3940] = 9'd4;
  assign mem[3941] = 9'd3;
  assign mem[3942] = 9'd4;
  assign mem[3943] = 9'd5;
  assign mem[3944] = 9'd7;
  assign mem[3945] = 9'd6;
  assign mem[3946] = 9'd5;
  assign mem[3947] = 9'd4;
  assign mem[3948] = 9'd3;
  assign mem[3949] = 9'd2;
  assign mem[3950] = 9'd3;
  assign mem[3951] = 9'd4;
  assign mem[3952] = 9'd6;
  assign mem[3953] = 9'd5;
  assign mem[3954] = 9'd4;
  assign mem[3955] = 9'd3;
  assign mem[3956] = 9'd2;
  assign mem[3957] = 9'd1;
  assign mem[3958] = 9'd2;
  assign mem[3959] = 9'd3;
  assign mem[3960] = 9'd5;
  assign mem[3961] = 9'd4;
  assign mem[3962] = 9'd3;
  assign mem[3963] = 9'd2;
  assign mem[3964] = 9'd1;
  assign mem[3965] = 9'd0;
  assign mem[3966] = 9'd1;
  assign mem[3967] = 9'd2;
  assign mem[3968] = 9'd13;
  assign mem[3969] = 9'd12;
  assign mem[3970] = 9'd11;
  assign mem[3971] = 9'd10;
  assign mem[3972] = 9'd9;
  assign mem[3973] = 9'd8;
  assign mem[3974] = 9'd7;
  assign mem[3975] = 9'd8;
  assign mem[3976] = 9'd12;
  assign mem[3977] = 9'd11;
  assign mem[3978] = 9'd10;
  assign mem[3979] = 9'd9;
  assign mem[3980] = 9'd8;
  assign mem[3981] = 9'd7;
  assign mem[3982] = 9'd6;
  assign mem[3983] = 9'd7;
  assign mem[3984] = 9'd11;
  assign mem[3985] = 9'd10;
  assign mem[3986] = 9'd9;
  assign mem[3987] = 9'd8;
  assign mem[3988] = 9'd7;
  assign mem[3989] = 9'd6;
  assign mem[3990] = 9'd5;
  assign mem[3991] = 9'd6;
  assign mem[3992] = 9'd10;
  assign mem[3993] = 9'd9;
  assign mem[3994] = 9'd8;
  assign mem[3995] = 9'd7;
  assign mem[3996] = 9'd6;
  assign mem[3997] = 9'd5;
  assign mem[3998] = 9'd4;
  assign mem[3999] = 9'd5;
  assign mem[4000] = 9'd9;
  assign mem[4001] = 9'd8;
  assign mem[4002] = 9'd7;
  assign mem[4003] = 9'd6;
  assign mem[4004] = 9'd5;
  assign mem[4005] = 9'd4;
  assign mem[4006] = 9'd3;
  assign mem[4007] = 9'd4;
  assign mem[4008] = 9'd8;
  assign mem[4009] = 9'd7;
  assign mem[4010] = 9'd6;
  assign mem[4011] = 9'd5;
  assign mem[4012] = 9'd4;
  assign mem[4013] = 9'd3;
  assign mem[4014] = 9'd2;
  assign mem[4015] = 9'd3;
  assign mem[4016] = 9'd7;
  assign mem[4017] = 9'd6;
  assign mem[4018] = 9'd5;
  assign mem[4019] = 9'd4;
  assign mem[4020] = 9'd3;
  assign mem[4021] = 9'd2;
  assign mem[4022] = 9'd1;
  assign mem[4023] = 9'd2;
  assign mem[4024] = 9'd6;
  assign mem[4025] = 9'd5;
  assign mem[4026] = 9'd4;
  assign mem[4027] = 9'd3;
  assign mem[4028] = 9'd2;
  assign mem[4029] = 9'd1;
  assign mem[4030] = 9'd0;
  assign mem[4031] = 9'd1;
  assign mem[4032] = 9'd14;
  assign mem[4033] = 9'd13;
  assign mem[4034] = 9'd12;
  assign mem[4035] = 9'd11;
  assign mem[4036] = 9'd10;
  assign mem[4037] = 9'd9;
  assign mem[4038] = 9'd8;
  assign mem[4039] = 9'd7;
  assign mem[4040] = 9'd13;
  assign mem[4041] = 9'd12;
  assign mem[4042] = 9'd11;
  assign mem[4043] = 9'd10;
  assign mem[4044] = 9'd9;
  assign mem[4045] = 9'd8;
  assign mem[4046] = 9'd7;
  assign mem[4047] = 9'd6;
  assign mem[4048] = 9'd12;
  assign mem[4049] = 9'd11;
  assign mem[4050] = 9'd10;
  assign mem[4051] = 9'd9;
  assign mem[4052] = 9'd8;
  assign mem[4053] = 9'd7;
  assign mem[4054] = 9'd6;
  assign mem[4055] = 9'd5;
  assign mem[4056] = 9'd11;
  assign mem[4057] = 9'd10;
  assign mem[4058] = 9'd9;
  assign mem[4059] = 9'd8;
  assign mem[4060] = 9'd7;
  assign mem[4061] = 9'd6;
  assign mem[4062] = 9'd5;
  assign mem[4063] = 9'd4;
  assign mem[4064] = 9'd10;
  assign mem[4065] = 9'd9;
  assign mem[4066] = 9'd8;
  assign mem[4067] = 9'd7;
  assign mem[4068] = 9'd6;
  assign mem[4069] = 9'd5;
  assign mem[4070] = 9'd4;
  assign mem[4071] = 9'd3;
  assign mem[4072] = 9'd9;
  assign mem[4073] = 9'd8;
  assign mem[4074] = 9'd7;
  assign mem[4075] = 9'd6;
  assign mem[4076] = 9'd5;
  assign mem[4077] = 9'd4;
  assign mem[4078] = 9'd3;
  assign mem[4079] = 9'd2;
  assign mem[4080] = 9'd8;
  assign mem[4081] = 9'd7;
  assign mem[4082] = 9'd6;
  assign mem[4083] = 9'd5;
  assign mem[4084] = 9'd4;
  assign mem[4085] = 9'd3;
  assign mem[4086] = 9'd2;
  assign mem[4087] = 9'd1;
  assign mem[4088] = 9'd7;
  assign mem[4089] = 9'd6;
  assign mem[4090] = 9'd5;
  assign mem[4091] = 9'd4;
  assign mem[4092] = 9'd3;
  assign mem[4093] = 9'd2;
  assign mem[4094] = 9'd1;
  assign mem[4095] = 9'd0;

endmodule



module st5_d2_s1_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [6-1:0] ca_in,
  input [6-1:0] cb_in,
  input [24-1:0] cva_in,
  input [4-1:0] cva_v_in,
  input [24-1:0] cvb_in,
  input [4-1:0] cvb_v_in,
  input [36-1:0] dvac_in,
  input [36-1:0] dvbc_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [18-1:0] dvac_out,
  output reg [18-1:0] dvbc_out,
  output reg [36-1:0] dvas_out,
  output reg [36-1:0] dvbs_out
);

  wire [6-1:0] cas;
  wire [6-1:0] cbs;
  wire [24-1:0] opva;
  wire [24-1:0] opvb;
  wire [18-1:0] dvac_t;
  wire [18-1:0] dvbc_t;
  wire [36-1:0] dvas_t;
  wire [36-1:0] dvbs_t;
  assign cas = cb_in;
  assign cbs = ca_in;
  assign dvac_t[8:0] = dvac_in[8:0] + dvac_in[17:9];
  assign dvac_t[17:9] = dvac_in[26:18] + dvac_in[35:27];
  assign dvbc_t[8:0] = dvbc_in[8:0] + dvbc_in[17:9];
  assign dvbc_t[17:9] = dvbc_in[26:18] + dvbc_in[35:27];
  assign opva[5:0] = (cva_in[5:0] == cas)? cbs : cva_in[5:0];
  assign opva[11:6] = (cva_in[11:6] == cas)? cbs : cva_in[11:6];
  assign opva[17:12] = (cva_in[17:12] == cas)? cbs : cva_in[17:12];
  assign opva[23:18] = (cva_in[23:18] == cas)? cbs : cva_in[23:18];
  assign opvb[5:0] = (cvb_in[5:0] == cbs)? cas : cvb_in[5:0];
  assign opvb[11:6] = (cvb_in[11:6] == cbs)? cas : cvb_in[11:6];
  assign opvb[17:12] = (cvb_in[17:12] == cbs)? cas : cvb_in[17:12];
  assign opvb[23:18] = (cvb_in[23:18] == cbs)? cas : cvb_in[23:18];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  distance_rom_8_8
  distance_rom_8_8_das_0
  (
    .opa0(cas),
    .opa1(opva[5:0]),
    .opav(cva_v_in[0]),
    .opb0(cas),
    .opb1(opva[11:6]),
    .opbv(cva_v_in[1]),
    .da(dvas_t[8:0]),
    .db(dvas_t[17:9])
  );


  distance_rom_8_8
  distance_rom_8_8_das_1
  (
    .opa0(cas),
    .opa1(opva[17:12]),
    .opav(cva_v_in[2]),
    .opb0(cas),
    .opb1(opva[23:18]),
    .opbv(cva_v_in[3]),
    .da(dvas_t[26:18]),
    .db(dvas_t[35:27])
  );


  distance_rom_8_8
  distance_rom_8_8_dbs_0
  (
    .opa0(cbs),
    .opa1(opvb[5:0]),
    .opav(cvb_v_in[0]),
    .opb0(cbs),
    .opb1(opvb[11:6]),
    .opbv(cvb_v_in[1]),
    .da(dvbs_t[8:0]),
    .db(dvbs_t[17:9])
  );


  distance_rom_8_8
  distance_rom_8_8_dbs_1
  (
    .opa0(cbs),
    .opa1(opvb[17:12]),
    .opav(cvb_v_in[2]),
    .opb0(cbs),
    .opb1(opvb[23:18]),
    .opbv(cvb_v_in[3]),
    .da(dvbs_t[26:18]),
    .db(dvbs_t[35:27])
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st6_s2_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [18-1:0] dvac_in,
  input [18-1:0] dvbc_in,
  input [36-1:0] dvas_in,
  input [36-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [9-1:0] dvac_out,
  output reg [9-1:0] dvbc_out,
  output reg [18-1:0] dvas_out,
  output reg [18-1:0] dvbs_out
);

  wire [9-1:0] dvac_t;
  wire [9-1:0] dvbc_t;
  wire [18-1:0] dvas_t;
  wire [18-1:0] dvbs_t;
  assign dvac_t = dvac_in[8:0] + dvac_in[17:9];
  assign dvbc_t = dvbc_in[8:0] + dvbc_in[17:9];
  assign dvas_t[8:0] = dvas_in[8:0] + dvas_in[17:9];
  assign dvas_t[17:9] = dvas_in[26:18] + dvas_in[35:27];
  assign dvbs_t[8:0] = dvbs_in[8:0] + dvbs_in[17:9];
  assign dvbs_t[17:9] = dvbs_in[26:18] + dvbs_in[35:27];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st7_s3_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [9-1:0] dvac_in,
  input [9-1:0] dvbc_in,
  input [18-1:0] dvas_in,
  input [18-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [9-1:0] dc_out,
  output reg [9-1:0] dvas_out,
  output reg [9-1:0] dvbs_out
);

  wire [9-1:0] dc_t;
  wire [9-1:0] dvas_t;
  wire [9-1:0] dvbs_t;
  assign dc_t = dvac_in + dvbc_in;
  assign dvas_t = dvas_in[8:0] + dvas_in[17:9];
  assign dvbs_t = dvbs_in[8:0] + dvbs_in[17:9];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dc_out <= dc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st8_s4_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [9-1:0] dc_in,
  input [9-1:0] dvas_in,
  input [9-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [9-1:0] dc_out,
  output reg [9-1:0] ds_out
);

  wire [9-1:0] ds_t;
  assign ds_t = dvas_in + dvbs_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dc_out <= dc_in;
    ds_out <= ds_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dc_out = 0;
    ds_out = 0;
  end


endmodule



module st9_cmp_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [9-1:0] dc_in,
  input [9-1:0] ds_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg sw_out
);

  wire sw_t;
  assign sw_t = ds_in < dc_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    sw_out <= sw_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    sw_out = 0;
  end


endmodule



module st10_reg_6th_64cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input sw_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg sw_out
);


  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    sw_out <= sw_in;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    sw_out = 0;
  end


endmodule

