

module sa_pipeline_6th_100cells
(
  input clk,
  input rst,
  input start,
  input [16-1:0] n_exec,
  output reg done
);

  // basic control inputs
  // -----
  wire pipe_start;
  reg [17-1:0] counter_total;
  // Threads controller output wires
  wire [3-1:0] th_idx;
  wire th_v;
  wire [7-1:0] th_ca;
  wire [7-1:0] th_cb;
  // -----

  always @(posedge clk) begin
    if(rst) begin
      counter_total <= 0;
      done <= 0;
    end else begin
      if((th_idx == 5) && ~th_v && &{ th_ca, th_cb }) begin
        counter_total <= counter_total + 1;
      end 
      if(counter_total == n_exec) begin
        done <= 1;
      end 
    end
  end

  // st1 output wires
  wire st1_rdy;
  wire [3-1:0] st1_idx;
  wire st1_v;
  wire [7-1:0] st1_ca;
  wire [7-1:0] st1_cb;
  wire [7-1:0] st1_na;
  wire st1_na_v;
  wire [7-1:0] st1_nb;
  wire st1_nb_v;
  wire st1_sw;
  wire [18-1:0] st1_wa;
  wire [18-1:0] st1_wb;
  // -----
  // st2 output wires
  wire [3-1:0] st2_idx;
  wire st2_v;
  wire [7-1:0] st2_ca;
  wire [7-1:0] st2_cb;
  wire [7-1:0] st2_na;
  wire st2_na_v;
  wire [7-1:0] st2_nb;
  wire st2_nb_v;
  wire [28-1:0] st2_va;
  wire [4-1:0] st2_va_v;
  wire [28-1:0] st2_vb;
  wire [4-1:0] st2_vb_v;
  wire st2_sw;
  wire [18-1:0] st2_wa;
  wire [18-1:0] st2_wb;
  // -----
  // st3 output wires
  wire [3-1:0] st3_idx;
  wire st3_v;
  wire [7-1:0] st3_ca;
  wire [7-1:0] st3_cb;
  wire [28-1:0] st3_cva;
  wire [4-1:0] st3_cva_v;
  wire [28-1:0] st3_cvb;
  wire [4-1:0] st3_cvb_v;
  wire [18-1:0] st3_wb;
  // -----
  // st4 output wires
  wire [3-1:0] st4_idx;
  wire st4_v;
  wire [7-1:0] st4_ca;
  wire [7-1:0] st4_cb;
  wire [28-1:0] st4_cva;
  wire [4-1:0] st4_cva_v;
  wire [28-1:0] st4_cvb;
  wire [4-1:0] st4_cvb_v;
  wire [40-1:0] st4_dvac;
  wire [40-1:0] st4_dvbc;
  // -----
  // st5 output wires
  wire [3-1:0] st5_idx;
  wire st5_v;
  wire [20-1:0] st5_dvac;
  wire [20-1:0] st5_dvbc;
  wire [40-1:0] st5_dvas;
  wire [40-1:0] st5_dvbs;
  // -----
  // st6 output wires
  wire [3-1:0] st6_idx;
  wire st6_v;
  wire [10-1:0] st6_dvac;
  wire [10-1:0] st6_dvbc;
  wire [20-1:0] st6_dvas;
  wire [20-1:0] st6_dvbs;
  // -----
  // st7 output wires
  wire [3-1:0] st7_idx;
  wire st7_v;
  wire [10-1:0] st7_dc;
  wire [10-1:0] st7_dvas;
  wire [10-1:0] st7_dvbs;
  // st8 output wires
  wire [3-1:0] st8_idx;
  wire st8_v;
  wire [10-1:0] st8_dc;
  wire [10-1:0] st8_ds;
  // -----
  // st9 output wires
  wire [3-1:0] st9_idx;
  wire st9_v;
  wire st9_sw;
  // -----
  // st10 output wires
  wire [3-1:0] st10_idx;
  wire st10_v;
  wire st10_sw;
  // -----
  assign pipe_start = &{ start, st1_rdy };

  th_controller_6th_100cells
  th_controller_6th_100cells
  (
    .clk(clk),
    .rst(rst),
    .start(pipe_start),
    .idx_out(th_idx),
    .v_out(th_v),
    .ca_out(th_ca),
    .cb_out(th_cb)
  );


  st1_c2n_6th_100cells
  st1_c2n_6th_100cells
  (
    .clk(clk),
    .rst(rst),
    .rdy(st1_rdy),
    .idx_in(th_idx),
    .v_in(th_v),
    .ca_in(th_ca),
    .cb_in(th_cb),
    .sw_in(st10_sw),
    .st1_wb_in(st1_wb),
    .idx_out(st1_idx),
    .v_out(st1_v),
    .ca_out(st1_ca),
    .cb_out(st1_cb),
    .na_out(st1_na),
    .na_v_out(st1_na_v),
    .nb_out(st1_nb),
    .nb_v_out(st1_nb_v),
    .sw_out(st1_sw),
    .wa_out(st1_wa),
    .wb_out(st1_wb)
  );


  st2_n_6th_100cells
  st2_n_6th_100cells
  (
    .clk(clk),
    .idx_in(st1_idx),
    .v_in(st1_v),
    .ca_in(st1_ca),
    .cb_in(st1_cb),
    .na_in(st1_na),
    .na_v_in(st1_na_v),
    .nb_in(st1_nb),
    .nb_v_in(st1_nb_v),
    .sw_in(st1_sw),
    .wa_in(st1_wa),
    .wb_in(st1_wb),
    .idx_out(st2_idx),
    .v_out(st2_v),
    .ca_out(st2_ca),
    .cb_out(st2_cb),
    .na_out(st2_na),
    .na_v_out(st2_na_v),
    .nb_out(st2_nb),
    .nb_v_out(st2_nb_v),
    .va_out(st2_va),
    .va_v_out(st2_va_v),
    .vb_out(st2_vb),
    .vb_v_out(st2_vb_v),
    .sw_out(st2_sw),
    .wa_out(st2_wa),
    .wb_out(st2_wb)
  );


  st3_n2c_6th_100cells
  st3_n2c_6th_100cells
  (
    .clk(clk),
    .rst(rst),
    .idx_in(st2_idx),
    .v_in(st2_v),
    .ca_in(st2_ca),
    .cb_in(st2_cb),
    .na_in(st2_na),
    .na_v_in(st2_na_v),
    .nb_in(st2_nb),
    .nb_v_in(st2_nb_v),
    .va_in(st2_va),
    .va_v_in(st2_va_v),
    .vb_in(st2_vb),
    .vb_v_in(st2_vb_v),
    .st3_wb_in(st3_wb),
    .sw_in(st2_sw),
    .wa_in(st2_wa),
    .wb_in(st2_wb),
    .idx_out(st3_idx),
    .v_out(st3_v),
    .ca_out(st3_ca),
    .cb_out(st3_cb),
    .cva_out(st3_cva),
    .cva_v_out(st3_cva_v),
    .cvb_out(st3_cvb),
    .cvb_v_out(st3_cvb_v),
    .wb_out(st3_wb)
  );


  st4_d1_6th_100cells
  st4_d1_6th_100cells
  (
    .clk(clk),
    .idx_in(st3_idx),
    .v_in(st3_v),
    .ca_in(st3_ca),
    .cb_in(st3_cb),
    .cva_in(st3_cva),
    .cva_v_in(st3_cva_v),
    .cvb_in(st3_cvb),
    .cvb_v_in(st3_cvb_v),
    .idx_out(st4_idx),
    .v_out(st4_v),
    .ca_out(st4_ca),
    .cb_out(st4_cb),
    .cva_out(st4_cva),
    .cva_v_out(st4_cva_v),
    .cvb_out(st4_cvb),
    .cvb_v_out(st4_cvb_v),
    .dvac_out(st4_dvac),
    .dvbc_out(st4_dvbc)
  );


  st5_d2_s1_6th_100cells
  st5_d2_s1_6th_100cells
  (
    .clk(clk),
    .idx_in(st4_idx),
    .v_in(st4_v),
    .ca_in(st4_ca),
    .cb_in(st4_cb),
    .cva_in(st4_cva),
    .cva_v_in(st4_cva_v),
    .cvb_in(st4_cvb),
    .cvb_v_in(st4_cvb_v),
    .dvac_in(st4_dvac),
    .dvbc_in(st4_dvbc),
    .idx_out(st5_idx),
    .v_out(st5_v),
    .dvac_out(st5_dvac),
    .dvbc_out(st5_dvbc),
    .dvas_out(st5_dvas),
    .dvbs_out(st5_dvbs)
  );


  st6_s2_6th_100cells
  st6_s2_6th_100cells
  (
    .clk(clk),
    .idx_in(st5_idx),
    .v_in(st5_v),
    .dvac_in(st5_dvac),
    .dvbc_in(st5_dvbc),
    .dvas_in(st5_dvas),
    .dvbs_in(st5_dvbs),
    .idx_out(st6_idx),
    .v_out(st6_v),
    .dvac_out(st6_dvac),
    .dvbc_out(st6_dvbc),
    .dvas_out(st6_dvas),
    .dvbs_out(st6_dvbs)
  );


  st7_s3_6th_100cells
  st7_s3_6th_100cells
  (
    .clk(clk),
    .idx_in(st6_idx),
    .v_in(st6_v),
    .dvac_in(st6_dvac),
    .dvbc_in(st6_dvbc),
    .dvas_in(st6_dvas),
    .dvbs_in(st6_dvbs),
    .idx_out(st7_idx),
    .v_out(st7_v),
    .dc_out(st7_dc),
    .dvas_out(st7_dvas),
    .dvbs_out(st7_dvbs)
  );


  st8_s4_6th_100cells
  st8_s4_6th_100cells
  (
    .clk(clk),
    .idx_in(st7_idx),
    .v_in(st7_v),
    .dc_in(st7_dc),
    .dvas_in(st7_dvas),
    .dvbs_in(st7_dvbs),
    .idx_out(st8_idx),
    .v_out(st8_v),
    .dc_out(st8_dc),
    .ds_out(st8_ds)
  );


  st9_cmp_6th_100cells
  st9_cmp_6th_100cells
  (
    .clk(clk),
    .idx_in(st8_idx),
    .v_in(st8_v),
    .dc_in(st8_dc),
    .ds_in(st8_ds),
    .idx_out(st9_idx),
    .v_out(st9_v),
    .sw_out(st9_sw)
  );


  st10_reg_6th_100cells
  st10_reg_6th_100cells
  (
    .clk(clk),
    .idx_in(st9_idx),
    .v_in(st9_v),
    .sw_in(st9_sw),
    .idx_out(st10_idx),
    .v_out(st10_v),
    .sw_out(st10_sw)
  );


  initial begin
    done = 0;
    counter_total = 0;
  end


endmodule



module th_controller_6th_100cells
(
  input clk,
  input rst,
  input start,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [7-1:0] ca_out,
  output reg [7-1:0] cb_out
);

  reg [6-1:0] flag_f_exec;
  reg [6-1:0] v_r;
  reg [3-1:0] idx_r;
  wire [14-1:0] counter;
  wire [14-1:0] counter_t;
  wire [14-1:0] counter_wr;
  wire [7-1:0] ca_out_t;
  wire [7-1:0] cb_out_t;
  assign counter_t = (flag_f_exec[idx_r])? 0 : counter;
  assign counter_wr = (&counter_t)? 0 : counter_t + 1;
  assign ca_out_t = counter_t[6:0];
  assign cb_out_t = counter_t[13:7];

  always @(posedge clk) begin
    if(rst) begin
      idx_out <= 0;
      v_out <= 0;
      ca_out <= 0;
      cb_out <= 0;
      idx_r <= 0;
      flag_f_exec <= 6'b111111;
      v_r <= 6'b111111;
    end else begin
      if(start) begin
        idx_out <= idx_r;
        v_out <= v_r[idx_r];
        ca_out <= ca_out_t;
        cb_out <= cb_out_t;
        v_r[idx_r] <= ~v_r[idx_r];
        if(!v_r[idx_r]) begin
          flag_f_exec[idx_r] <= 0;
          if(idx_r == 5) begin
            idx_r <= 0;
          end else begin
            idx_r <= idx_r + 1;
          end
        end 
      end 
    end
  end


  mem_2r_1w_width14_depth3
  #(
    .init_file("./rom/th.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width14_depth3
  (
    .clk(clk),
    .rd_addr0(idx_r),
    .out0(counter),
    .wr(~v_r[idx_r]),
    .wr_addr(idx_r),
    .wr_data(counter_wr)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    flag_f_exec = 0;
    v_r = 0;
    idx_r = 0;
  end


endmodule



module mem_2r_1w_width14_depth3 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [3-1:0] rd_addr0,
  input [3-1:0] rd_addr1,
  output [14-1:0] out0,
  output [14-1:0] out1,
  input wr,
  input [3-1:0] wr_addr,
  input [14-1:0] wr_data
);

  reg [14-1:0] mem [0:2**3-1];
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end


  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end

  //synthesis translate_on

endmodule



module st1_c2n_6th_100cells
(
  input clk,
  input rst,
  input [3-1:0] idx_in,
  input v_in,
  input [7-1:0] ca_in,
  input [7-1:0] cb_in,
  input sw_in,
  input [18-1:0] st1_wb_in,
  output reg rdy,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [7-1:0] ca_out,
  output reg [7-1:0] cb_out,
  output reg [7-1:0] na_out,
  output reg na_v_out,
  output reg [7-1:0] nb_out,
  output reg nb_v_out,
  output reg sw_out,
  output reg [18-1:0] wa_out,
  output reg [18-1:0] wb_out
);

  reg flag;
  reg [4-1:0] counter;
  reg fifo_init;
  wire [7-1:0] na_t;
  wire na_v_t;
  wire [7-1:0] nb_t;
  wire nb_v_t;
  wire [18-1:0] wa_t;
  wire [18-1:0] wb_t;
  wire fifoa_wr_en;
  wire fifoa_rd_en;
  wire [18-1:0] fifoa_data;
  wire fifob_wr_en;
  wire fifob_rd_en;
  wire [18-1:0] fifob_data;
  wire [3-1:0] wa_idx;
  wire [7-1:0] wa_c;
  wire [7-1:0] wa_n;
  wire wa_n_v;
  wire [3-1:0] wb_idx;
  wire [7-1:0] wb_c;
  wire [7-1:0] wb_n;
  wire wb_n_v;
  wire m_wr;
  wire [10-1:0] m_wr_addr;
  wire [8-1:0] m_wr_data;
  assign fifoa_data = { idx_in, ca_in, nb_v_t, nb_t };
  assign fifob_data = { idx_in, cb_in, na_v_t, na_t };
  assign fifoa_rd_en = &{ rdy, v_in };
  assign fifob_rd_en = &{ rdy, v_in };
  assign fifoa_wr_en = |{ &{ rdy, v_in }, fifo_init };
  assign fifob_wr_en = |{ &{ rdy, v_in }, fifo_init };
  assign wa_n = wa_t[6:0];
  assign wa_n_v = wa_t[7];
  assign wa_c = wa_t[14:8];
  assign wa_idx = wa_t[17:15];
  assign wb_n = st1_wb_in[6:0];
  assign wb_n_v = st1_wb_in[7];
  assign wb_c = st1_wb_in[14:8];
  assign wb_idx = st1_wb_in[17:15];
  assign m_wr = sw_in;
  assign m_wr_addr = (flag)? { wa_idx, wa_c } : { wb_idx, wb_c };
  assign m_wr_data = (flag)? { wa_n_v, wa_n } : { wb_n_v, wb_n };

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    na_out <= na_t;
    na_v_out <= na_v_t;
    nb_out <= nb_t;
    nb_v_out <= nb_v_t;
    sw_out <= sw_in;
    wa_out <= wa_t;
    wb_out <= wb_t;
  end


  always @(posedge clk) begin
    if(rst) begin
      flag <= 1;
    end else begin
      if(sw_in) begin
        flag <= ~flag;
      end 
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      rdy <= 0;
      fifo_init <= 0;
      counter <= 0;
    end else begin
      if(counter == 4) begin
        rdy <= 1;
        fifo_init <= 0;
      end else begin
        counter <= counter + 1;
        fifo_init <= 1;
      end
    end
  end


  mem_2r_1w_width8_depth10
  #(
    .init_file("./rom/c_n.rom"),
    .read_f(1),
    .write_f(1),
    .output_file("./rom/c_n_out.rom")
  )
  mem_2r_1w_width8_depth10
  (
    .clk(clk),
    .rd_addr0({ idx_in, ca_in }),
    .rd_addr1({ idx_in, cb_in }),
    .out0({ na_v_t, na_t }),
    .out1({ nb_v_t, nb_t }),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  fifo
  #(
    .FIFO_WIDTH(18),
    .FIFO_DEPTH_BITS(3)
  )
  fifo_a
  (
    .clk(clk),
    .rst(rst),
    .write_enable(fifoa_wr_en),
    .input_data(fifoa_data),
    .output_read_enable(fifoa_rd_en),
    .output_data(wa_t)
  );


  fifo
  #(
    .FIFO_WIDTH(18),
    .FIFO_DEPTH_BITS(3)
  )
  fifo_b
  (
    .clk(clk),
    .rst(rst),
    .write_enable(fifob_wr_en),
    .input_data(fifob_data),
    .output_read_enable(fifob_rd_en),
    .output_data(wb_t)
  );


  initial begin
    rdy = 0;
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    na_out = 0;
    na_v_out = 0;
    nb_out = 0;
    nb_v_out = 0;
    sw_out = 0;
    wa_out = 0;
    wb_out = 0;
    flag = 0;
    counter = 0;
    fifo_init = 0;
  end


endmodule



module mem_2r_1w_width8_depth10 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [10-1:0] rd_addr0,
  input [10-1:0] rd_addr1,
  output [8-1:0] out0,
  output [8-1:0] out1,
  input wr,
  input [10-1:0] wr_addr,
  input [8-1:0] wr_data
);

  reg [8-1:0] mem [0:2**10-1];
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end


  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end

  //synthesis translate_on

endmodule



module fifo #
(
  parameter FIFO_WIDTH = 32,
  parameter FIFO_DEPTH_BITS = 8,
  parameter FIFO_ALMOSTFULL_THRESHOLD = 2 ** FIFO_DEPTH_BITS - 4,
  parameter FIFO_ALMOSTEMPTY_THRESHOLD = 4
)
(
  input clk,
  input rst,
  input write_enable,
  input [FIFO_WIDTH-1:0] input_data,
  input output_read_enable,
  output reg output_valid,
  output reg [FIFO_WIDTH-1:0] output_data,
  output reg empty,
  output reg almostempty,
  output reg full,
  output reg almostfull,
  output reg [FIFO_DEPTH_BITS+1-1:0] data_count
);

  reg [FIFO_DEPTH_BITS-1:0] read_pointer;
  reg [FIFO_DEPTH_BITS-1:0] write_pointer;
  reg [FIFO_WIDTH-1:0] mem [0:2**FIFO_DEPTH_BITS-1];

  always @(posedge clk) begin
    if(rst) begin
      empty <= 1;
      almostempty <= 1;
      full <= 0;
      almostfull <= 0;
      read_pointer <= 0;
      write_pointer <= 0;
      data_count <= 0;
    end else begin
      case({ write_enable, output_read_enable })
        3: begin
          read_pointer <= read_pointer + 1;
          write_pointer <= write_pointer + 1;
        end
        2: begin
          if(~full) begin
            write_pointer <= write_pointer + 1;
            data_count <= data_count + 1;
            empty <= 0;
            if(data_count == FIFO_ALMOSTEMPTY_THRESHOLD - 1) begin
              almostempty <= 0;
            end 
            if(data_count == 2 ** FIFO_DEPTH_BITS - 1) begin
              full <= 1;
            end 
            if(data_count == FIFO_ALMOSTFULL_THRESHOLD - 1) begin
              almostfull <= 1;
            end 
          end 
        end
        1: begin
          if(~empty) begin
            read_pointer <= read_pointer + 1;
            data_count <= data_count - 1;
            full <= 0;
            if(data_count == FIFO_ALMOSTFULL_THRESHOLD) begin
              almostfull <= 0;
            end 
            if(data_count == 1) begin
              empty <= 1;
            end 
            if(data_count == FIFO_ALMOSTEMPTY_THRESHOLD) begin
              almostempty <= 1;
            end 
          end 
        end
      endcase
    end
  end


  always @(posedge clk) begin
    if(rst) begin
      output_valid <= 0;
    end else begin
      output_valid <= 0;
      if(write_enable == 1) begin
        mem[write_pointer] <= input_data;
      end 
      if(output_read_enable == 1) begin
        output_data <= mem[read_pointer];
        output_valid <= 1;
      end 
    end
  end


endmodule



module st2_n_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [7-1:0] ca_in,
  input [7-1:0] cb_in,
  input [7-1:0] na_in,
  input na_v_in,
  input [7-1:0] nb_in,
  input nb_v_in,
  input sw_in,
  input [18-1:0] wa_in,
  input [18-1:0] wb_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [7-1:0] ca_out,
  output reg [7-1:0] cb_out,
  output reg [7-1:0] na_out,
  output reg na_v_out,
  output reg [7-1:0] nb_out,
  output reg nb_v_out,
  output reg [28-1:0] va_out,
  output reg [4-1:0] va_v_out,
  output reg [28-1:0] vb_out,
  output reg [4-1:0] vb_v_out,
  output reg sw_out,
  output reg [18-1:0] wa_out,
  output reg [18-1:0] wb_out
);

  wire [28-1:0] va_t;
  wire [4-1:0] va_v_t;
  wire [4-1:0] va_v_m;
  wire [28-1:0] vb_t;
  wire [4-1:0] vb_v_t;
  wire [4-1:0] vb_v_m;
  assign va_v_t = (na_v_in)? va_v_m : 4'b0;
  assign vb_v_t = (nb_v_in)? vb_v_m : 4'b0;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    na_out <= na_in;
    na_v_out <= na_v_in;
    nb_out <= nb_in;
    nb_v_out <= nb_v_in;
    sw_out <= sw_in;
    wa_out <= wa_in;
    wb_out <= wb_in;
    va_out <= va_t;
    va_v_out <= va_v_t;
    vb_out <= vb_t;
    vb_v_out <= vb_v_t;
  end


  mem_2r_1w_width8_depth7
  #(
    .init_file("./rom/n0.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width8_depth7_0
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[0], va_t[6:0] }),
    .out1({ vb_v_m[0], vb_t[6:0] }),
    .wr(1'b0),
    .wr_addr(7'b0),
    .wr_data(8'b0)
  );


  mem_2r_1w_width8_depth7
  #(
    .init_file("./rom/n1.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width8_depth7_1
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[1], va_t[13:7] }),
    .out1({ vb_v_m[1], vb_t[13:7] }),
    .wr(1'b0),
    .wr_addr(7'b0),
    .wr_data(8'b0)
  );


  mem_2r_1w_width8_depth7
  #(
    .init_file("./rom/n2.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width8_depth7_2
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[2], va_t[20:14] }),
    .out1({ vb_v_m[2], vb_t[20:14] }),
    .wr(1'b0),
    .wr_addr(7'b0),
    .wr_data(8'b0)
  );


  mem_2r_1w_width8_depth7
  #(
    .init_file("./rom/n3.rom"),
    .read_f(1),
    .write_f(0)
  )
  mem_2r_1w_width8_depth7_3
  (
    .clk(clk),
    .rd_addr0(na_in),
    .rd_addr1(nb_in),
    .out0({ va_v_m[3], va_t[27:21] }),
    .out1({ vb_v_m[3], vb_t[27:21] }),
    .wr(1'b0),
    .wr_addr(7'b0),
    .wr_data(8'b0)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    na_out = 0;
    na_v_out = 0;
    nb_out = 0;
    nb_v_out = 0;
    va_out = 0;
    va_v_out = 0;
    vb_out = 0;
    vb_v_out = 0;
    sw_out = 0;
    wa_out = 0;
    wb_out = 0;
  end


endmodule



module mem_2r_1w_width8_depth7 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [7-1:0] rd_addr0,
  input [7-1:0] rd_addr1,
  output [8-1:0] out0,
  output [8-1:0] out1,
  input wr,
  input [7-1:0] wr_addr,
  input [8-1:0] wr_data
);

  reg [8-1:0] mem [0:2**7-1];
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end


  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end

  //synthesis translate_on

endmodule



module st3_n2c_6th_100cells
(
  input clk,
  input rst,
  input [3-1:0] idx_in,
  input v_in,
  input [7-1:0] ca_in,
  input [7-1:0] cb_in,
  input [7-1:0] na_in,
  input na_v_in,
  input [7-1:0] nb_in,
  input nb_v_in,
  input [28-1:0] va_in,
  input [4-1:0] va_v_in,
  input [28-1:0] vb_in,
  input [4-1:0] vb_v_in,
  input [18-1:0] st3_wb_in,
  input sw_in,
  input [18-1:0] wa_in,
  input [18-1:0] wb_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [7-1:0] ca_out,
  output reg [7-1:0] cb_out,
  output reg [28-1:0] cva_out,
  output reg [4-1:0] cva_v_out,
  output reg [28-1:0] cvb_out,
  output reg [4-1:0] cvb_v_out,
  output reg [18-1:0] wb_out
);

  reg flag;
  wire [28-1:0] cva_t;
  wire [28-1:0] cvb_t;
  wire [3-1:0] wa_idx;
  wire [7-1:0] wa_c;
  wire [7-1:0] wa_n;
  wire wa_n_v;
  wire [3-1:0] wb_idx;
  wire [7-1:0] wb_c;
  wire [7-1:0] wb_n;
  wire wb_n_v;
  wire m_wr;
  wire [10-1:0] m_wr_addr;
  wire [7-1:0] m_wr_data;
  assign wa_n = wa_in[6:0];
  assign wa_n_v = wa_in[7];
  assign wa_c = wa_in[14:8];
  assign wa_idx = wa_in[17:15];
  assign wb_n = st3_wb_in[6:0];
  assign wb_n_v = st3_wb_in[7];
  assign wb_c = st3_wb_in[14:8];
  assign wb_idx = st3_wb_in[17:15];
  assign m_wr = (flag)? &{ sw_in, wa_n_v } : &{ sw_in, wb_n_v };
  assign m_wr_addr = (flag)? { wa_idx, wa_n } : { wb_idx, wb_n };
  assign m_wr_data = (flag)? wa_c : wb_c;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    cva_out <= cva_t;
    cva_v_out <= va_v_in;
    cvb_out <= cvb_t;
    cvb_v_out <= vb_v_in;
    wb_out <= wb_in;
  end


  always @(posedge clk) begin
    if(rst) begin
      flag <= 1;
    end else begin
      if(sw_in) begin
        flag <= ~flag;
      end 
    end
  end


  mem_2r_1w_width7_depth10
  #(
    .init_file("./rom/n_c.rom"),
    .read_f(1),
    .write_f(1),
    .output_file("./rom/n_c_out.rom")
  )
  mem_2r_1w_width7_depth10_0
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[6:0] }),
    .rd_addr1({ idx_in, vb_in[6:0] }),
    .out0(cva_t[6:0]),
    .out1(cvb_t[6:0]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width7_depth10
  #(
    .init_file("./rom/n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./rom/n_c_out.rom")
  )
  mem_2r_1w_width7_depth10_1
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[13:7] }),
    .rd_addr1({ idx_in, vb_in[13:7] }),
    .out0(cva_t[13:7]),
    .out1(cvb_t[13:7]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width7_depth10
  #(
    .init_file("./rom/n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./rom/n_c_out.rom")
  )
  mem_2r_1w_width7_depth10_2
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[20:14] }),
    .rd_addr1({ idx_in, vb_in[20:14] }),
    .out0(cva_t[20:14]),
    .out1(cvb_t[20:14]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  mem_2r_1w_width7_depth10
  #(
    .init_file("./rom/n_c.rom"),
    .read_f(1),
    .write_f(0),
    .output_file("./rom/n_c_out.rom")
  )
  mem_2r_1w_width7_depth10_3
  (
    .clk(clk),
    .rd_addr0({ idx_in, va_in[27:21] }),
    .rd_addr1({ idx_in, vb_in[27:21] }),
    .out0(cva_t[27:21]),
    .out1(cvb_t[27:21]),
    .wr(m_wr),
    .wr_addr(m_wr_addr),
    .wr_data(m_wr_data)
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    cva_out = 0;
    cva_v_out = 0;
    cvb_out = 0;
    cvb_v_out = 0;
    wb_out = 0;
    flag = 0;
  end


endmodule



module mem_2r_1w_width7_depth10 #
(
  parameter read_f = 0,
  parameter init_file = "mem_file.txt",
  parameter write_f = 0,
  parameter output_file = "mem_out_file.txt"
)
(
  input clk,
  input [10-1:0] rd_addr0,
  input [10-1:0] rd_addr1,
  output [7-1:0] out0,
  output [7-1:0] out1,
  input wr,
  input [10-1:0] wr_addr,
  input [7-1:0] wr_data
);

  reg [7-1:0] mem [0:2**10-1];
  assign out0 = mem[rd_addr0];
  assign out1 = mem[rd_addr1];

  always @(posedge clk) begin
    if(wr) begin
      mem[wr_addr] <= wr_data;
    end 
  end

  //synthesis translate_off

  always @(posedge clk) begin
    if(wr && write_f) begin
      $writememh(output_file, mem);
    end 
  end


  initial begin
    if(read_f) begin
      $readmemh(init_file, mem);
    end 
  end

  //synthesis translate_on

endmodule



module st4_d1_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [7-1:0] ca_in,
  input [7-1:0] cb_in,
  input [28-1:0] cva_in,
  input [4-1:0] cva_v_in,
  input [28-1:0] cvb_in,
  input [4-1:0] cvb_v_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [7-1:0] ca_out,
  output reg [7-1:0] cb_out,
  output reg [28-1:0] cva_out,
  output reg [4-1:0] cva_v_out,
  output reg [28-1:0] cvb_out,
  output reg [4-1:0] cvb_v_out,
  output reg [40-1:0] dvac_out,
  output reg [40-1:0] dvbc_out
);

  wire [7-1:0] cac;
  wire [7-1:0] cbc;
  wire [40-1:0] dvac_t;
  wire [40-1:0] dvbc_t;
  assign cac = ca_in;
  assign cbc = cb_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    ca_out <= ca_in;
    cb_out <= cb_in;
    cva_out <= cva_in;
    cva_v_out <= cva_v_in;
    cvb_out <= cvb_in;
    cvb_v_out <= cvb_v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
  end


  distance_rom_10_10
  distance_rom_10_10_dac_0
  (
    .opa0(cac),
    .opa1(cva_in[6:0]),
    .opav(cva_v_in[0]),
    .opb0(cac),
    .opb1(cva_in[13:7]),
    .opbv(cva_v_in[1]),
    .da(dvac_t[9:0]),
    .db(dvac_t[19:10])
  );


  distance_rom_10_10
  distance_rom_10_10_dac_1
  (
    .opa0(cac),
    .opa1(cva_in[20:14]),
    .opav(cva_v_in[2]),
    .opb0(cac),
    .opb1(cva_in[27:21]),
    .opbv(cva_v_in[3]),
    .da(dvac_t[29:20]),
    .db(dvac_t[39:30])
  );


  distance_rom_10_10
  distance_rom_10_10_dbc_0
  (
    .opa0(cbc),
    .opa1(cvb_in[6:0]),
    .opav(cvb_v_in[0]),
    .opb0(cbc),
    .opb1(cvb_in[13:7]),
    .opbv(cvb_v_in[1]),
    .da(dvbc_t[9:0]),
    .db(dvbc_t[19:10])
  );


  distance_rom_10_10
  distance_rom_10_10_dbc_1
  (
    .opa0(cbc),
    .opa1(cvb_in[20:14]),
    .opav(cvb_v_in[2]),
    .opb0(cbc),
    .opb1(cvb_in[27:21]),
    .opbv(cvb_v_in[3]),
    .da(dvbc_t[29:20]),
    .db(dvbc_t[39:30])
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    ca_out = 0;
    cb_out = 0;
    cva_out = 0;
    cva_v_out = 0;
    cvb_out = 0;
    cvb_v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
  end


endmodule



module distance_rom_10_10
(
  input [7-1:0] opa0,
  input [7-1:0] opa1,
  input opav,
  input [7-1:0] opb0,
  input [7-1:0] opb1,
  input opbv,
  output [10-1:0] da,
  output [10-1:0] db
);

  wire [10-1:0] mem [0:100**2-1];
  assign da = (opav)? mem[{ opa1, opa0 }] : 0;
  assign db = (opbv)? mem[{ opb1, opb0 }] : 0;
  assign mem[0] = 10'd0;
  assign mem[1] = 10'd1;
  assign mem[2] = 10'd2;
  assign mem[3] = 10'd3;
  assign mem[4] = 10'd4;
  assign mem[5] = 10'd5;
  assign mem[6] = 10'd6;
  assign mem[7] = 10'd7;
  assign mem[8] = 10'd8;
  assign mem[9] = 10'd9;
  assign mem[10] = 10'd1;
  assign mem[11] = 10'd2;
  assign mem[12] = 10'd3;
  assign mem[13] = 10'd4;
  assign mem[14] = 10'd5;
  assign mem[15] = 10'd6;
  assign mem[16] = 10'd7;
  assign mem[17] = 10'd8;
  assign mem[18] = 10'd9;
  assign mem[19] = 10'd10;
  assign mem[20] = 10'd2;
  assign mem[21] = 10'd3;
  assign mem[22] = 10'd4;
  assign mem[23] = 10'd5;
  assign mem[24] = 10'd6;
  assign mem[25] = 10'd7;
  assign mem[26] = 10'd8;
  assign mem[27] = 10'd9;
  assign mem[28] = 10'd10;
  assign mem[29] = 10'd11;
  assign mem[30] = 10'd3;
  assign mem[31] = 10'd4;
  assign mem[32] = 10'd5;
  assign mem[33] = 10'd6;
  assign mem[34] = 10'd7;
  assign mem[35] = 10'd8;
  assign mem[36] = 10'd9;
  assign mem[37] = 10'd10;
  assign mem[38] = 10'd11;
  assign mem[39] = 10'd12;
  assign mem[40] = 10'd4;
  assign mem[41] = 10'd5;
  assign mem[42] = 10'd6;
  assign mem[43] = 10'd7;
  assign mem[44] = 10'd8;
  assign mem[45] = 10'd9;
  assign mem[46] = 10'd10;
  assign mem[47] = 10'd11;
  assign mem[48] = 10'd12;
  assign mem[49] = 10'd13;
  assign mem[50] = 10'd5;
  assign mem[51] = 10'd6;
  assign mem[52] = 10'd7;
  assign mem[53] = 10'd8;
  assign mem[54] = 10'd9;
  assign mem[55] = 10'd10;
  assign mem[56] = 10'd11;
  assign mem[57] = 10'd12;
  assign mem[58] = 10'd13;
  assign mem[59] = 10'd14;
  assign mem[60] = 10'd6;
  assign mem[61] = 10'd7;
  assign mem[62] = 10'd8;
  assign mem[63] = 10'd9;
  assign mem[64] = 10'd10;
  assign mem[65] = 10'd11;
  assign mem[66] = 10'd12;
  assign mem[67] = 10'd13;
  assign mem[68] = 10'd14;
  assign mem[69] = 10'd15;
  assign mem[70] = 10'd7;
  assign mem[71] = 10'd8;
  assign mem[72] = 10'd9;
  assign mem[73] = 10'd10;
  assign mem[74] = 10'd11;
  assign mem[75] = 10'd12;
  assign mem[76] = 10'd13;
  assign mem[77] = 10'd14;
  assign mem[78] = 10'd15;
  assign mem[79] = 10'd16;
  assign mem[80] = 10'd8;
  assign mem[81] = 10'd9;
  assign mem[82] = 10'd10;
  assign mem[83] = 10'd11;
  assign mem[84] = 10'd12;
  assign mem[85] = 10'd13;
  assign mem[86] = 10'd14;
  assign mem[87] = 10'd15;
  assign mem[88] = 10'd16;
  assign mem[89] = 10'd17;
  assign mem[90] = 10'd9;
  assign mem[91] = 10'd10;
  assign mem[92] = 10'd11;
  assign mem[93] = 10'd12;
  assign mem[94] = 10'd13;
  assign mem[95] = 10'd14;
  assign mem[96] = 10'd15;
  assign mem[97] = 10'd16;
  assign mem[98] = 10'd17;
  assign mem[99] = 10'd18;
  assign mem[100] = 10'd1;
  assign mem[101] = 10'd0;
  assign mem[102] = 10'd1;
  assign mem[103] = 10'd2;
  assign mem[104] = 10'd3;
  assign mem[105] = 10'd4;
  assign mem[106] = 10'd5;
  assign mem[107] = 10'd6;
  assign mem[108] = 10'd7;
  assign mem[109] = 10'd8;
  assign mem[110] = 10'd2;
  assign mem[111] = 10'd1;
  assign mem[112] = 10'd2;
  assign mem[113] = 10'd3;
  assign mem[114] = 10'd4;
  assign mem[115] = 10'd5;
  assign mem[116] = 10'd6;
  assign mem[117] = 10'd7;
  assign mem[118] = 10'd8;
  assign mem[119] = 10'd9;
  assign mem[120] = 10'd3;
  assign mem[121] = 10'd2;
  assign mem[122] = 10'd3;
  assign mem[123] = 10'd4;
  assign mem[124] = 10'd5;
  assign mem[125] = 10'd6;
  assign mem[126] = 10'd7;
  assign mem[127] = 10'd8;
  assign mem[128] = 10'd9;
  assign mem[129] = 10'd10;
  assign mem[130] = 10'd4;
  assign mem[131] = 10'd3;
  assign mem[132] = 10'd4;
  assign mem[133] = 10'd5;
  assign mem[134] = 10'd6;
  assign mem[135] = 10'd7;
  assign mem[136] = 10'd8;
  assign mem[137] = 10'd9;
  assign mem[138] = 10'd10;
  assign mem[139] = 10'd11;
  assign mem[140] = 10'd5;
  assign mem[141] = 10'd4;
  assign mem[142] = 10'd5;
  assign mem[143] = 10'd6;
  assign mem[144] = 10'd7;
  assign mem[145] = 10'd8;
  assign mem[146] = 10'd9;
  assign mem[147] = 10'd10;
  assign mem[148] = 10'd11;
  assign mem[149] = 10'd12;
  assign mem[150] = 10'd6;
  assign mem[151] = 10'd5;
  assign mem[152] = 10'd6;
  assign mem[153] = 10'd7;
  assign mem[154] = 10'd8;
  assign mem[155] = 10'd9;
  assign mem[156] = 10'd10;
  assign mem[157] = 10'd11;
  assign mem[158] = 10'd12;
  assign mem[159] = 10'd13;
  assign mem[160] = 10'd7;
  assign mem[161] = 10'd6;
  assign mem[162] = 10'd7;
  assign mem[163] = 10'd8;
  assign mem[164] = 10'd9;
  assign mem[165] = 10'd10;
  assign mem[166] = 10'd11;
  assign mem[167] = 10'd12;
  assign mem[168] = 10'd13;
  assign mem[169] = 10'd14;
  assign mem[170] = 10'd8;
  assign mem[171] = 10'd7;
  assign mem[172] = 10'd8;
  assign mem[173] = 10'd9;
  assign mem[174] = 10'd10;
  assign mem[175] = 10'd11;
  assign mem[176] = 10'd12;
  assign mem[177] = 10'd13;
  assign mem[178] = 10'd14;
  assign mem[179] = 10'd15;
  assign mem[180] = 10'd9;
  assign mem[181] = 10'd8;
  assign mem[182] = 10'd9;
  assign mem[183] = 10'd10;
  assign mem[184] = 10'd11;
  assign mem[185] = 10'd12;
  assign mem[186] = 10'd13;
  assign mem[187] = 10'd14;
  assign mem[188] = 10'd15;
  assign mem[189] = 10'd16;
  assign mem[190] = 10'd10;
  assign mem[191] = 10'd9;
  assign mem[192] = 10'd10;
  assign mem[193] = 10'd11;
  assign mem[194] = 10'd12;
  assign mem[195] = 10'd13;
  assign mem[196] = 10'd14;
  assign mem[197] = 10'd15;
  assign mem[198] = 10'd16;
  assign mem[199] = 10'd17;
  assign mem[200] = 10'd2;
  assign mem[201] = 10'd1;
  assign mem[202] = 10'd0;
  assign mem[203] = 10'd1;
  assign mem[204] = 10'd2;
  assign mem[205] = 10'd3;
  assign mem[206] = 10'd4;
  assign mem[207] = 10'd5;
  assign mem[208] = 10'd6;
  assign mem[209] = 10'd7;
  assign mem[210] = 10'd3;
  assign mem[211] = 10'd2;
  assign mem[212] = 10'd1;
  assign mem[213] = 10'd2;
  assign mem[214] = 10'd3;
  assign mem[215] = 10'd4;
  assign mem[216] = 10'd5;
  assign mem[217] = 10'd6;
  assign mem[218] = 10'd7;
  assign mem[219] = 10'd8;
  assign mem[220] = 10'd4;
  assign mem[221] = 10'd3;
  assign mem[222] = 10'd2;
  assign mem[223] = 10'd3;
  assign mem[224] = 10'd4;
  assign mem[225] = 10'd5;
  assign mem[226] = 10'd6;
  assign mem[227] = 10'd7;
  assign mem[228] = 10'd8;
  assign mem[229] = 10'd9;
  assign mem[230] = 10'd5;
  assign mem[231] = 10'd4;
  assign mem[232] = 10'd3;
  assign mem[233] = 10'd4;
  assign mem[234] = 10'd5;
  assign mem[235] = 10'd6;
  assign mem[236] = 10'd7;
  assign mem[237] = 10'd8;
  assign mem[238] = 10'd9;
  assign mem[239] = 10'd10;
  assign mem[240] = 10'd6;
  assign mem[241] = 10'd5;
  assign mem[242] = 10'd4;
  assign mem[243] = 10'd5;
  assign mem[244] = 10'd6;
  assign mem[245] = 10'd7;
  assign mem[246] = 10'd8;
  assign mem[247] = 10'd9;
  assign mem[248] = 10'd10;
  assign mem[249] = 10'd11;
  assign mem[250] = 10'd7;
  assign mem[251] = 10'd6;
  assign mem[252] = 10'd5;
  assign mem[253] = 10'd6;
  assign mem[254] = 10'd7;
  assign mem[255] = 10'd8;
  assign mem[256] = 10'd9;
  assign mem[257] = 10'd10;
  assign mem[258] = 10'd11;
  assign mem[259] = 10'd12;
  assign mem[260] = 10'd8;
  assign mem[261] = 10'd7;
  assign mem[262] = 10'd6;
  assign mem[263] = 10'd7;
  assign mem[264] = 10'd8;
  assign mem[265] = 10'd9;
  assign mem[266] = 10'd10;
  assign mem[267] = 10'd11;
  assign mem[268] = 10'd12;
  assign mem[269] = 10'd13;
  assign mem[270] = 10'd9;
  assign mem[271] = 10'd8;
  assign mem[272] = 10'd7;
  assign mem[273] = 10'd8;
  assign mem[274] = 10'd9;
  assign mem[275] = 10'd10;
  assign mem[276] = 10'd11;
  assign mem[277] = 10'd12;
  assign mem[278] = 10'd13;
  assign mem[279] = 10'd14;
  assign mem[280] = 10'd10;
  assign mem[281] = 10'd9;
  assign mem[282] = 10'd8;
  assign mem[283] = 10'd9;
  assign mem[284] = 10'd10;
  assign mem[285] = 10'd11;
  assign mem[286] = 10'd12;
  assign mem[287] = 10'd13;
  assign mem[288] = 10'd14;
  assign mem[289] = 10'd15;
  assign mem[290] = 10'd11;
  assign mem[291] = 10'd10;
  assign mem[292] = 10'd9;
  assign mem[293] = 10'd10;
  assign mem[294] = 10'd11;
  assign mem[295] = 10'd12;
  assign mem[296] = 10'd13;
  assign mem[297] = 10'd14;
  assign mem[298] = 10'd15;
  assign mem[299] = 10'd16;
  assign mem[300] = 10'd3;
  assign mem[301] = 10'd2;
  assign mem[302] = 10'd1;
  assign mem[303] = 10'd0;
  assign mem[304] = 10'd1;
  assign mem[305] = 10'd2;
  assign mem[306] = 10'd3;
  assign mem[307] = 10'd4;
  assign mem[308] = 10'd5;
  assign mem[309] = 10'd6;
  assign mem[310] = 10'd4;
  assign mem[311] = 10'd3;
  assign mem[312] = 10'd2;
  assign mem[313] = 10'd1;
  assign mem[314] = 10'd2;
  assign mem[315] = 10'd3;
  assign mem[316] = 10'd4;
  assign mem[317] = 10'd5;
  assign mem[318] = 10'd6;
  assign mem[319] = 10'd7;
  assign mem[320] = 10'd5;
  assign mem[321] = 10'd4;
  assign mem[322] = 10'd3;
  assign mem[323] = 10'd2;
  assign mem[324] = 10'd3;
  assign mem[325] = 10'd4;
  assign mem[326] = 10'd5;
  assign mem[327] = 10'd6;
  assign mem[328] = 10'd7;
  assign mem[329] = 10'd8;
  assign mem[330] = 10'd6;
  assign mem[331] = 10'd5;
  assign mem[332] = 10'd4;
  assign mem[333] = 10'd3;
  assign mem[334] = 10'd4;
  assign mem[335] = 10'd5;
  assign mem[336] = 10'd6;
  assign mem[337] = 10'd7;
  assign mem[338] = 10'd8;
  assign mem[339] = 10'd9;
  assign mem[340] = 10'd7;
  assign mem[341] = 10'd6;
  assign mem[342] = 10'd5;
  assign mem[343] = 10'd4;
  assign mem[344] = 10'd5;
  assign mem[345] = 10'd6;
  assign mem[346] = 10'd7;
  assign mem[347] = 10'd8;
  assign mem[348] = 10'd9;
  assign mem[349] = 10'd10;
  assign mem[350] = 10'd8;
  assign mem[351] = 10'd7;
  assign mem[352] = 10'd6;
  assign mem[353] = 10'd5;
  assign mem[354] = 10'd6;
  assign mem[355] = 10'd7;
  assign mem[356] = 10'd8;
  assign mem[357] = 10'd9;
  assign mem[358] = 10'd10;
  assign mem[359] = 10'd11;
  assign mem[360] = 10'd9;
  assign mem[361] = 10'd8;
  assign mem[362] = 10'd7;
  assign mem[363] = 10'd6;
  assign mem[364] = 10'd7;
  assign mem[365] = 10'd8;
  assign mem[366] = 10'd9;
  assign mem[367] = 10'd10;
  assign mem[368] = 10'd11;
  assign mem[369] = 10'd12;
  assign mem[370] = 10'd10;
  assign mem[371] = 10'd9;
  assign mem[372] = 10'd8;
  assign mem[373] = 10'd7;
  assign mem[374] = 10'd8;
  assign mem[375] = 10'd9;
  assign mem[376] = 10'd10;
  assign mem[377] = 10'd11;
  assign mem[378] = 10'd12;
  assign mem[379] = 10'd13;
  assign mem[380] = 10'd11;
  assign mem[381] = 10'd10;
  assign mem[382] = 10'd9;
  assign mem[383] = 10'd8;
  assign mem[384] = 10'd9;
  assign mem[385] = 10'd10;
  assign mem[386] = 10'd11;
  assign mem[387] = 10'd12;
  assign mem[388] = 10'd13;
  assign mem[389] = 10'd14;
  assign mem[390] = 10'd12;
  assign mem[391] = 10'd11;
  assign mem[392] = 10'd10;
  assign mem[393] = 10'd9;
  assign mem[394] = 10'd10;
  assign mem[395] = 10'd11;
  assign mem[396] = 10'd12;
  assign mem[397] = 10'd13;
  assign mem[398] = 10'd14;
  assign mem[399] = 10'd15;
  assign mem[400] = 10'd4;
  assign mem[401] = 10'd3;
  assign mem[402] = 10'd2;
  assign mem[403] = 10'd1;
  assign mem[404] = 10'd0;
  assign mem[405] = 10'd1;
  assign mem[406] = 10'd2;
  assign mem[407] = 10'd3;
  assign mem[408] = 10'd4;
  assign mem[409] = 10'd5;
  assign mem[410] = 10'd5;
  assign mem[411] = 10'd4;
  assign mem[412] = 10'd3;
  assign mem[413] = 10'd2;
  assign mem[414] = 10'd1;
  assign mem[415] = 10'd2;
  assign mem[416] = 10'd3;
  assign mem[417] = 10'd4;
  assign mem[418] = 10'd5;
  assign mem[419] = 10'd6;
  assign mem[420] = 10'd6;
  assign mem[421] = 10'd5;
  assign mem[422] = 10'd4;
  assign mem[423] = 10'd3;
  assign mem[424] = 10'd2;
  assign mem[425] = 10'd3;
  assign mem[426] = 10'd4;
  assign mem[427] = 10'd5;
  assign mem[428] = 10'd6;
  assign mem[429] = 10'd7;
  assign mem[430] = 10'd7;
  assign mem[431] = 10'd6;
  assign mem[432] = 10'd5;
  assign mem[433] = 10'd4;
  assign mem[434] = 10'd3;
  assign mem[435] = 10'd4;
  assign mem[436] = 10'd5;
  assign mem[437] = 10'd6;
  assign mem[438] = 10'd7;
  assign mem[439] = 10'd8;
  assign mem[440] = 10'd8;
  assign mem[441] = 10'd7;
  assign mem[442] = 10'd6;
  assign mem[443] = 10'd5;
  assign mem[444] = 10'd4;
  assign mem[445] = 10'd5;
  assign mem[446] = 10'd6;
  assign mem[447] = 10'd7;
  assign mem[448] = 10'd8;
  assign mem[449] = 10'd9;
  assign mem[450] = 10'd9;
  assign mem[451] = 10'd8;
  assign mem[452] = 10'd7;
  assign mem[453] = 10'd6;
  assign mem[454] = 10'd5;
  assign mem[455] = 10'd6;
  assign mem[456] = 10'd7;
  assign mem[457] = 10'd8;
  assign mem[458] = 10'd9;
  assign mem[459] = 10'd10;
  assign mem[460] = 10'd10;
  assign mem[461] = 10'd9;
  assign mem[462] = 10'd8;
  assign mem[463] = 10'd7;
  assign mem[464] = 10'd6;
  assign mem[465] = 10'd7;
  assign mem[466] = 10'd8;
  assign mem[467] = 10'd9;
  assign mem[468] = 10'd10;
  assign mem[469] = 10'd11;
  assign mem[470] = 10'd11;
  assign mem[471] = 10'd10;
  assign mem[472] = 10'd9;
  assign mem[473] = 10'd8;
  assign mem[474] = 10'd7;
  assign mem[475] = 10'd8;
  assign mem[476] = 10'd9;
  assign mem[477] = 10'd10;
  assign mem[478] = 10'd11;
  assign mem[479] = 10'd12;
  assign mem[480] = 10'd12;
  assign mem[481] = 10'd11;
  assign mem[482] = 10'd10;
  assign mem[483] = 10'd9;
  assign mem[484] = 10'd8;
  assign mem[485] = 10'd9;
  assign mem[486] = 10'd10;
  assign mem[487] = 10'd11;
  assign mem[488] = 10'd12;
  assign mem[489] = 10'd13;
  assign mem[490] = 10'd13;
  assign mem[491] = 10'd12;
  assign mem[492] = 10'd11;
  assign mem[493] = 10'd10;
  assign mem[494] = 10'd9;
  assign mem[495] = 10'd10;
  assign mem[496] = 10'd11;
  assign mem[497] = 10'd12;
  assign mem[498] = 10'd13;
  assign mem[499] = 10'd14;
  assign mem[500] = 10'd5;
  assign mem[501] = 10'd4;
  assign mem[502] = 10'd3;
  assign mem[503] = 10'd2;
  assign mem[504] = 10'd1;
  assign mem[505] = 10'd0;
  assign mem[506] = 10'd1;
  assign mem[507] = 10'd2;
  assign mem[508] = 10'd3;
  assign mem[509] = 10'd4;
  assign mem[510] = 10'd6;
  assign mem[511] = 10'd5;
  assign mem[512] = 10'd4;
  assign mem[513] = 10'd3;
  assign mem[514] = 10'd2;
  assign mem[515] = 10'd1;
  assign mem[516] = 10'd2;
  assign mem[517] = 10'd3;
  assign mem[518] = 10'd4;
  assign mem[519] = 10'd5;
  assign mem[520] = 10'd7;
  assign mem[521] = 10'd6;
  assign mem[522] = 10'd5;
  assign mem[523] = 10'd4;
  assign mem[524] = 10'd3;
  assign mem[525] = 10'd2;
  assign mem[526] = 10'd3;
  assign mem[527] = 10'd4;
  assign mem[528] = 10'd5;
  assign mem[529] = 10'd6;
  assign mem[530] = 10'd8;
  assign mem[531] = 10'd7;
  assign mem[532] = 10'd6;
  assign mem[533] = 10'd5;
  assign mem[534] = 10'd4;
  assign mem[535] = 10'd3;
  assign mem[536] = 10'd4;
  assign mem[537] = 10'd5;
  assign mem[538] = 10'd6;
  assign mem[539] = 10'd7;
  assign mem[540] = 10'd9;
  assign mem[541] = 10'd8;
  assign mem[542] = 10'd7;
  assign mem[543] = 10'd6;
  assign mem[544] = 10'd5;
  assign mem[545] = 10'd4;
  assign mem[546] = 10'd5;
  assign mem[547] = 10'd6;
  assign mem[548] = 10'd7;
  assign mem[549] = 10'd8;
  assign mem[550] = 10'd10;
  assign mem[551] = 10'd9;
  assign mem[552] = 10'd8;
  assign mem[553] = 10'd7;
  assign mem[554] = 10'd6;
  assign mem[555] = 10'd5;
  assign mem[556] = 10'd6;
  assign mem[557] = 10'd7;
  assign mem[558] = 10'd8;
  assign mem[559] = 10'd9;
  assign mem[560] = 10'd11;
  assign mem[561] = 10'd10;
  assign mem[562] = 10'd9;
  assign mem[563] = 10'd8;
  assign mem[564] = 10'd7;
  assign mem[565] = 10'd6;
  assign mem[566] = 10'd7;
  assign mem[567] = 10'd8;
  assign mem[568] = 10'd9;
  assign mem[569] = 10'd10;
  assign mem[570] = 10'd12;
  assign mem[571] = 10'd11;
  assign mem[572] = 10'd10;
  assign mem[573] = 10'd9;
  assign mem[574] = 10'd8;
  assign mem[575] = 10'd7;
  assign mem[576] = 10'd8;
  assign mem[577] = 10'd9;
  assign mem[578] = 10'd10;
  assign mem[579] = 10'd11;
  assign mem[580] = 10'd13;
  assign mem[581] = 10'd12;
  assign mem[582] = 10'd11;
  assign mem[583] = 10'd10;
  assign mem[584] = 10'd9;
  assign mem[585] = 10'd8;
  assign mem[586] = 10'd9;
  assign mem[587] = 10'd10;
  assign mem[588] = 10'd11;
  assign mem[589] = 10'd12;
  assign mem[590] = 10'd14;
  assign mem[591] = 10'd13;
  assign mem[592] = 10'd12;
  assign mem[593] = 10'd11;
  assign mem[594] = 10'd10;
  assign mem[595] = 10'd9;
  assign mem[596] = 10'd10;
  assign mem[597] = 10'd11;
  assign mem[598] = 10'd12;
  assign mem[599] = 10'd13;
  assign mem[600] = 10'd6;
  assign mem[601] = 10'd5;
  assign mem[602] = 10'd4;
  assign mem[603] = 10'd3;
  assign mem[604] = 10'd2;
  assign mem[605] = 10'd1;
  assign mem[606] = 10'd0;
  assign mem[607] = 10'd1;
  assign mem[608] = 10'd2;
  assign mem[609] = 10'd3;
  assign mem[610] = 10'd7;
  assign mem[611] = 10'd6;
  assign mem[612] = 10'd5;
  assign mem[613] = 10'd4;
  assign mem[614] = 10'd3;
  assign mem[615] = 10'd2;
  assign mem[616] = 10'd1;
  assign mem[617] = 10'd2;
  assign mem[618] = 10'd3;
  assign mem[619] = 10'd4;
  assign mem[620] = 10'd8;
  assign mem[621] = 10'd7;
  assign mem[622] = 10'd6;
  assign mem[623] = 10'd5;
  assign mem[624] = 10'd4;
  assign mem[625] = 10'd3;
  assign mem[626] = 10'd2;
  assign mem[627] = 10'd3;
  assign mem[628] = 10'd4;
  assign mem[629] = 10'd5;
  assign mem[630] = 10'd9;
  assign mem[631] = 10'd8;
  assign mem[632] = 10'd7;
  assign mem[633] = 10'd6;
  assign mem[634] = 10'd5;
  assign mem[635] = 10'd4;
  assign mem[636] = 10'd3;
  assign mem[637] = 10'd4;
  assign mem[638] = 10'd5;
  assign mem[639] = 10'd6;
  assign mem[640] = 10'd10;
  assign mem[641] = 10'd9;
  assign mem[642] = 10'd8;
  assign mem[643] = 10'd7;
  assign mem[644] = 10'd6;
  assign mem[645] = 10'd5;
  assign mem[646] = 10'd4;
  assign mem[647] = 10'd5;
  assign mem[648] = 10'd6;
  assign mem[649] = 10'd7;
  assign mem[650] = 10'd11;
  assign mem[651] = 10'd10;
  assign mem[652] = 10'd9;
  assign mem[653] = 10'd8;
  assign mem[654] = 10'd7;
  assign mem[655] = 10'd6;
  assign mem[656] = 10'd5;
  assign mem[657] = 10'd6;
  assign mem[658] = 10'd7;
  assign mem[659] = 10'd8;
  assign mem[660] = 10'd12;
  assign mem[661] = 10'd11;
  assign mem[662] = 10'd10;
  assign mem[663] = 10'd9;
  assign mem[664] = 10'd8;
  assign mem[665] = 10'd7;
  assign mem[666] = 10'd6;
  assign mem[667] = 10'd7;
  assign mem[668] = 10'd8;
  assign mem[669] = 10'd9;
  assign mem[670] = 10'd13;
  assign mem[671] = 10'd12;
  assign mem[672] = 10'd11;
  assign mem[673] = 10'd10;
  assign mem[674] = 10'd9;
  assign mem[675] = 10'd8;
  assign mem[676] = 10'd7;
  assign mem[677] = 10'd8;
  assign mem[678] = 10'd9;
  assign mem[679] = 10'd10;
  assign mem[680] = 10'd14;
  assign mem[681] = 10'd13;
  assign mem[682] = 10'd12;
  assign mem[683] = 10'd11;
  assign mem[684] = 10'd10;
  assign mem[685] = 10'd9;
  assign mem[686] = 10'd8;
  assign mem[687] = 10'd9;
  assign mem[688] = 10'd10;
  assign mem[689] = 10'd11;
  assign mem[690] = 10'd15;
  assign mem[691] = 10'd14;
  assign mem[692] = 10'd13;
  assign mem[693] = 10'd12;
  assign mem[694] = 10'd11;
  assign mem[695] = 10'd10;
  assign mem[696] = 10'd9;
  assign mem[697] = 10'd10;
  assign mem[698] = 10'd11;
  assign mem[699] = 10'd12;
  assign mem[700] = 10'd7;
  assign mem[701] = 10'd6;
  assign mem[702] = 10'd5;
  assign mem[703] = 10'd4;
  assign mem[704] = 10'd3;
  assign mem[705] = 10'd2;
  assign mem[706] = 10'd1;
  assign mem[707] = 10'd0;
  assign mem[708] = 10'd1;
  assign mem[709] = 10'd2;
  assign mem[710] = 10'd8;
  assign mem[711] = 10'd7;
  assign mem[712] = 10'd6;
  assign mem[713] = 10'd5;
  assign mem[714] = 10'd4;
  assign mem[715] = 10'd3;
  assign mem[716] = 10'd2;
  assign mem[717] = 10'd1;
  assign mem[718] = 10'd2;
  assign mem[719] = 10'd3;
  assign mem[720] = 10'd9;
  assign mem[721] = 10'd8;
  assign mem[722] = 10'd7;
  assign mem[723] = 10'd6;
  assign mem[724] = 10'd5;
  assign mem[725] = 10'd4;
  assign mem[726] = 10'd3;
  assign mem[727] = 10'd2;
  assign mem[728] = 10'd3;
  assign mem[729] = 10'd4;
  assign mem[730] = 10'd10;
  assign mem[731] = 10'd9;
  assign mem[732] = 10'd8;
  assign mem[733] = 10'd7;
  assign mem[734] = 10'd6;
  assign mem[735] = 10'd5;
  assign mem[736] = 10'd4;
  assign mem[737] = 10'd3;
  assign mem[738] = 10'd4;
  assign mem[739] = 10'd5;
  assign mem[740] = 10'd11;
  assign mem[741] = 10'd10;
  assign mem[742] = 10'd9;
  assign mem[743] = 10'd8;
  assign mem[744] = 10'd7;
  assign mem[745] = 10'd6;
  assign mem[746] = 10'd5;
  assign mem[747] = 10'd4;
  assign mem[748] = 10'd5;
  assign mem[749] = 10'd6;
  assign mem[750] = 10'd12;
  assign mem[751] = 10'd11;
  assign mem[752] = 10'd10;
  assign mem[753] = 10'd9;
  assign mem[754] = 10'd8;
  assign mem[755] = 10'd7;
  assign mem[756] = 10'd6;
  assign mem[757] = 10'd5;
  assign mem[758] = 10'd6;
  assign mem[759] = 10'd7;
  assign mem[760] = 10'd13;
  assign mem[761] = 10'd12;
  assign mem[762] = 10'd11;
  assign mem[763] = 10'd10;
  assign mem[764] = 10'd9;
  assign mem[765] = 10'd8;
  assign mem[766] = 10'd7;
  assign mem[767] = 10'd6;
  assign mem[768] = 10'd7;
  assign mem[769] = 10'd8;
  assign mem[770] = 10'd14;
  assign mem[771] = 10'd13;
  assign mem[772] = 10'd12;
  assign mem[773] = 10'd11;
  assign mem[774] = 10'd10;
  assign mem[775] = 10'd9;
  assign mem[776] = 10'd8;
  assign mem[777] = 10'd7;
  assign mem[778] = 10'd8;
  assign mem[779] = 10'd9;
  assign mem[780] = 10'd15;
  assign mem[781] = 10'd14;
  assign mem[782] = 10'd13;
  assign mem[783] = 10'd12;
  assign mem[784] = 10'd11;
  assign mem[785] = 10'd10;
  assign mem[786] = 10'd9;
  assign mem[787] = 10'd8;
  assign mem[788] = 10'd9;
  assign mem[789] = 10'd10;
  assign mem[790] = 10'd16;
  assign mem[791] = 10'd15;
  assign mem[792] = 10'd14;
  assign mem[793] = 10'd13;
  assign mem[794] = 10'd12;
  assign mem[795] = 10'd11;
  assign mem[796] = 10'd10;
  assign mem[797] = 10'd9;
  assign mem[798] = 10'd10;
  assign mem[799] = 10'd11;
  assign mem[800] = 10'd8;
  assign mem[801] = 10'd7;
  assign mem[802] = 10'd6;
  assign mem[803] = 10'd5;
  assign mem[804] = 10'd4;
  assign mem[805] = 10'd3;
  assign mem[806] = 10'd2;
  assign mem[807] = 10'd1;
  assign mem[808] = 10'd0;
  assign mem[809] = 10'd1;
  assign mem[810] = 10'd9;
  assign mem[811] = 10'd8;
  assign mem[812] = 10'd7;
  assign mem[813] = 10'd6;
  assign mem[814] = 10'd5;
  assign mem[815] = 10'd4;
  assign mem[816] = 10'd3;
  assign mem[817] = 10'd2;
  assign mem[818] = 10'd1;
  assign mem[819] = 10'd2;
  assign mem[820] = 10'd10;
  assign mem[821] = 10'd9;
  assign mem[822] = 10'd8;
  assign mem[823] = 10'd7;
  assign mem[824] = 10'd6;
  assign mem[825] = 10'd5;
  assign mem[826] = 10'd4;
  assign mem[827] = 10'd3;
  assign mem[828] = 10'd2;
  assign mem[829] = 10'd3;
  assign mem[830] = 10'd11;
  assign mem[831] = 10'd10;
  assign mem[832] = 10'd9;
  assign mem[833] = 10'd8;
  assign mem[834] = 10'd7;
  assign mem[835] = 10'd6;
  assign mem[836] = 10'd5;
  assign mem[837] = 10'd4;
  assign mem[838] = 10'd3;
  assign mem[839] = 10'd4;
  assign mem[840] = 10'd12;
  assign mem[841] = 10'd11;
  assign mem[842] = 10'd10;
  assign mem[843] = 10'd9;
  assign mem[844] = 10'd8;
  assign mem[845] = 10'd7;
  assign mem[846] = 10'd6;
  assign mem[847] = 10'd5;
  assign mem[848] = 10'd4;
  assign mem[849] = 10'd5;
  assign mem[850] = 10'd13;
  assign mem[851] = 10'd12;
  assign mem[852] = 10'd11;
  assign mem[853] = 10'd10;
  assign mem[854] = 10'd9;
  assign mem[855] = 10'd8;
  assign mem[856] = 10'd7;
  assign mem[857] = 10'd6;
  assign mem[858] = 10'd5;
  assign mem[859] = 10'd6;
  assign mem[860] = 10'd14;
  assign mem[861] = 10'd13;
  assign mem[862] = 10'd12;
  assign mem[863] = 10'd11;
  assign mem[864] = 10'd10;
  assign mem[865] = 10'd9;
  assign mem[866] = 10'd8;
  assign mem[867] = 10'd7;
  assign mem[868] = 10'd6;
  assign mem[869] = 10'd7;
  assign mem[870] = 10'd15;
  assign mem[871] = 10'd14;
  assign mem[872] = 10'd13;
  assign mem[873] = 10'd12;
  assign mem[874] = 10'd11;
  assign mem[875] = 10'd10;
  assign mem[876] = 10'd9;
  assign mem[877] = 10'd8;
  assign mem[878] = 10'd7;
  assign mem[879] = 10'd8;
  assign mem[880] = 10'd16;
  assign mem[881] = 10'd15;
  assign mem[882] = 10'd14;
  assign mem[883] = 10'd13;
  assign mem[884] = 10'd12;
  assign mem[885] = 10'd11;
  assign mem[886] = 10'd10;
  assign mem[887] = 10'd9;
  assign mem[888] = 10'd8;
  assign mem[889] = 10'd9;
  assign mem[890] = 10'd17;
  assign mem[891] = 10'd16;
  assign mem[892] = 10'd15;
  assign mem[893] = 10'd14;
  assign mem[894] = 10'd13;
  assign mem[895] = 10'd12;
  assign mem[896] = 10'd11;
  assign mem[897] = 10'd10;
  assign mem[898] = 10'd9;
  assign mem[899] = 10'd10;
  assign mem[900] = 10'd9;
  assign mem[901] = 10'd8;
  assign mem[902] = 10'd7;
  assign mem[903] = 10'd6;
  assign mem[904] = 10'd5;
  assign mem[905] = 10'd4;
  assign mem[906] = 10'd3;
  assign mem[907] = 10'd2;
  assign mem[908] = 10'd1;
  assign mem[909] = 10'd0;
  assign mem[910] = 10'd10;
  assign mem[911] = 10'd9;
  assign mem[912] = 10'd8;
  assign mem[913] = 10'd7;
  assign mem[914] = 10'd6;
  assign mem[915] = 10'd5;
  assign mem[916] = 10'd4;
  assign mem[917] = 10'd3;
  assign mem[918] = 10'd2;
  assign mem[919] = 10'd1;
  assign mem[920] = 10'd11;
  assign mem[921] = 10'd10;
  assign mem[922] = 10'd9;
  assign mem[923] = 10'd8;
  assign mem[924] = 10'd7;
  assign mem[925] = 10'd6;
  assign mem[926] = 10'd5;
  assign mem[927] = 10'd4;
  assign mem[928] = 10'd3;
  assign mem[929] = 10'd2;
  assign mem[930] = 10'd12;
  assign mem[931] = 10'd11;
  assign mem[932] = 10'd10;
  assign mem[933] = 10'd9;
  assign mem[934] = 10'd8;
  assign mem[935] = 10'd7;
  assign mem[936] = 10'd6;
  assign mem[937] = 10'd5;
  assign mem[938] = 10'd4;
  assign mem[939] = 10'd3;
  assign mem[940] = 10'd13;
  assign mem[941] = 10'd12;
  assign mem[942] = 10'd11;
  assign mem[943] = 10'd10;
  assign mem[944] = 10'd9;
  assign mem[945] = 10'd8;
  assign mem[946] = 10'd7;
  assign mem[947] = 10'd6;
  assign mem[948] = 10'd5;
  assign mem[949] = 10'd4;
  assign mem[950] = 10'd14;
  assign mem[951] = 10'd13;
  assign mem[952] = 10'd12;
  assign mem[953] = 10'd11;
  assign mem[954] = 10'd10;
  assign mem[955] = 10'd9;
  assign mem[956] = 10'd8;
  assign mem[957] = 10'd7;
  assign mem[958] = 10'd6;
  assign mem[959] = 10'd5;
  assign mem[960] = 10'd15;
  assign mem[961] = 10'd14;
  assign mem[962] = 10'd13;
  assign mem[963] = 10'd12;
  assign mem[964] = 10'd11;
  assign mem[965] = 10'd10;
  assign mem[966] = 10'd9;
  assign mem[967] = 10'd8;
  assign mem[968] = 10'd7;
  assign mem[969] = 10'd6;
  assign mem[970] = 10'd16;
  assign mem[971] = 10'd15;
  assign mem[972] = 10'd14;
  assign mem[973] = 10'd13;
  assign mem[974] = 10'd12;
  assign mem[975] = 10'd11;
  assign mem[976] = 10'd10;
  assign mem[977] = 10'd9;
  assign mem[978] = 10'd8;
  assign mem[979] = 10'd7;
  assign mem[980] = 10'd17;
  assign mem[981] = 10'd16;
  assign mem[982] = 10'd15;
  assign mem[983] = 10'd14;
  assign mem[984] = 10'd13;
  assign mem[985] = 10'd12;
  assign mem[986] = 10'd11;
  assign mem[987] = 10'd10;
  assign mem[988] = 10'd9;
  assign mem[989] = 10'd8;
  assign mem[990] = 10'd18;
  assign mem[991] = 10'd17;
  assign mem[992] = 10'd16;
  assign mem[993] = 10'd15;
  assign mem[994] = 10'd14;
  assign mem[995] = 10'd13;
  assign mem[996] = 10'd12;
  assign mem[997] = 10'd11;
  assign mem[998] = 10'd10;
  assign mem[999] = 10'd9;
  assign mem[1000] = 10'd1;
  assign mem[1001] = 10'd2;
  assign mem[1002] = 10'd3;
  assign mem[1003] = 10'd4;
  assign mem[1004] = 10'd5;
  assign mem[1005] = 10'd6;
  assign mem[1006] = 10'd7;
  assign mem[1007] = 10'd8;
  assign mem[1008] = 10'd9;
  assign mem[1009] = 10'd10;
  assign mem[1010] = 10'd0;
  assign mem[1011] = 10'd1;
  assign mem[1012] = 10'd2;
  assign mem[1013] = 10'd3;
  assign mem[1014] = 10'd4;
  assign mem[1015] = 10'd5;
  assign mem[1016] = 10'd6;
  assign mem[1017] = 10'd7;
  assign mem[1018] = 10'd8;
  assign mem[1019] = 10'd9;
  assign mem[1020] = 10'd1;
  assign mem[1021] = 10'd2;
  assign mem[1022] = 10'd3;
  assign mem[1023] = 10'd4;
  assign mem[1024] = 10'd5;
  assign mem[1025] = 10'd6;
  assign mem[1026] = 10'd7;
  assign mem[1027] = 10'd8;
  assign mem[1028] = 10'd9;
  assign mem[1029] = 10'd10;
  assign mem[1030] = 10'd2;
  assign mem[1031] = 10'd3;
  assign mem[1032] = 10'd4;
  assign mem[1033] = 10'd5;
  assign mem[1034] = 10'd6;
  assign mem[1035] = 10'd7;
  assign mem[1036] = 10'd8;
  assign mem[1037] = 10'd9;
  assign mem[1038] = 10'd10;
  assign mem[1039] = 10'd11;
  assign mem[1040] = 10'd3;
  assign mem[1041] = 10'd4;
  assign mem[1042] = 10'd5;
  assign mem[1043] = 10'd6;
  assign mem[1044] = 10'd7;
  assign mem[1045] = 10'd8;
  assign mem[1046] = 10'd9;
  assign mem[1047] = 10'd10;
  assign mem[1048] = 10'd11;
  assign mem[1049] = 10'd12;
  assign mem[1050] = 10'd4;
  assign mem[1051] = 10'd5;
  assign mem[1052] = 10'd6;
  assign mem[1053] = 10'd7;
  assign mem[1054] = 10'd8;
  assign mem[1055] = 10'd9;
  assign mem[1056] = 10'd10;
  assign mem[1057] = 10'd11;
  assign mem[1058] = 10'd12;
  assign mem[1059] = 10'd13;
  assign mem[1060] = 10'd5;
  assign mem[1061] = 10'd6;
  assign mem[1062] = 10'd7;
  assign mem[1063] = 10'd8;
  assign mem[1064] = 10'd9;
  assign mem[1065] = 10'd10;
  assign mem[1066] = 10'd11;
  assign mem[1067] = 10'd12;
  assign mem[1068] = 10'd13;
  assign mem[1069] = 10'd14;
  assign mem[1070] = 10'd6;
  assign mem[1071] = 10'd7;
  assign mem[1072] = 10'd8;
  assign mem[1073] = 10'd9;
  assign mem[1074] = 10'd10;
  assign mem[1075] = 10'd11;
  assign mem[1076] = 10'd12;
  assign mem[1077] = 10'd13;
  assign mem[1078] = 10'd14;
  assign mem[1079] = 10'd15;
  assign mem[1080] = 10'd7;
  assign mem[1081] = 10'd8;
  assign mem[1082] = 10'd9;
  assign mem[1083] = 10'd10;
  assign mem[1084] = 10'd11;
  assign mem[1085] = 10'd12;
  assign mem[1086] = 10'd13;
  assign mem[1087] = 10'd14;
  assign mem[1088] = 10'd15;
  assign mem[1089] = 10'd16;
  assign mem[1090] = 10'd8;
  assign mem[1091] = 10'd9;
  assign mem[1092] = 10'd10;
  assign mem[1093] = 10'd11;
  assign mem[1094] = 10'd12;
  assign mem[1095] = 10'd13;
  assign mem[1096] = 10'd14;
  assign mem[1097] = 10'd15;
  assign mem[1098] = 10'd16;
  assign mem[1099] = 10'd17;
  assign mem[1100] = 10'd2;
  assign mem[1101] = 10'd1;
  assign mem[1102] = 10'd2;
  assign mem[1103] = 10'd3;
  assign mem[1104] = 10'd4;
  assign mem[1105] = 10'd5;
  assign mem[1106] = 10'd6;
  assign mem[1107] = 10'd7;
  assign mem[1108] = 10'd8;
  assign mem[1109] = 10'd9;
  assign mem[1110] = 10'd1;
  assign mem[1111] = 10'd0;
  assign mem[1112] = 10'd1;
  assign mem[1113] = 10'd2;
  assign mem[1114] = 10'd3;
  assign mem[1115] = 10'd4;
  assign mem[1116] = 10'd5;
  assign mem[1117] = 10'd6;
  assign mem[1118] = 10'd7;
  assign mem[1119] = 10'd8;
  assign mem[1120] = 10'd2;
  assign mem[1121] = 10'd1;
  assign mem[1122] = 10'd2;
  assign mem[1123] = 10'd3;
  assign mem[1124] = 10'd4;
  assign mem[1125] = 10'd5;
  assign mem[1126] = 10'd6;
  assign mem[1127] = 10'd7;
  assign mem[1128] = 10'd8;
  assign mem[1129] = 10'd9;
  assign mem[1130] = 10'd3;
  assign mem[1131] = 10'd2;
  assign mem[1132] = 10'd3;
  assign mem[1133] = 10'd4;
  assign mem[1134] = 10'd5;
  assign mem[1135] = 10'd6;
  assign mem[1136] = 10'd7;
  assign mem[1137] = 10'd8;
  assign mem[1138] = 10'd9;
  assign mem[1139] = 10'd10;
  assign mem[1140] = 10'd4;
  assign mem[1141] = 10'd3;
  assign mem[1142] = 10'd4;
  assign mem[1143] = 10'd5;
  assign mem[1144] = 10'd6;
  assign mem[1145] = 10'd7;
  assign mem[1146] = 10'd8;
  assign mem[1147] = 10'd9;
  assign mem[1148] = 10'd10;
  assign mem[1149] = 10'd11;
  assign mem[1150] = 10'd5;
  assign mem[1151] = 10'd4;
  assign mem[1152] = 10'd5;
  assign mem[1153] = 10'd6;
  assign mem[1154] = 10'd7;
  assign mem[1155] = 10'd8;
  assign mem[1156] = 10'd9;
  assign mem[1157] = 10'd10;
  assign mem[1158] = 10'd11;
  assign mem[1159] = 10'd12;
  assign mem[1160] = 10'd6;
  assign mem[1161] = 10'd5;
  assign mem[1162] = 10'd6;
  assign mem[1163] = 10'd7;
  assign mem[1164] = 10'd8;
  assign mem[1165] = 10'd9;
  assign mem[1166] = 10'd10;
  assign mem[1167] = 10'd11;
  assign mem[1168] = 10'd12;
  assign mem[1169] = 10'd13;
  assign mem[1170] = 10'd7;
  assign mem[1171] = 10'd6;
  assign mem[1172] = 10'd7;
  assign mem[1173] = 10'd8;
  assign mem[1174] = 10'd9;
  assign mem[1175] = 10'd10;
  assign mem[1176] = 10'd11;
  assign mem[1177] = 10'd12;
  assign mem[1178] = 10'd13;
  assign mem[1179] = 10'd14;
  assign mem[1180] = 10'd8;
  assign mem[1181] = 10'd7;
  assign mem[1182] = 10'd8;
  assign mem[1183] = 10'd9;
  assign mem[1184] = 10'd10;
  assign mem[1185] = 10'd11;
  assign mem[1186] = 10'd12;
  assign mem[1187] = 10'd13;
  assign mem[1188] = 10'd14;
  assign mem[1189] = 10'd15;
  assign mem[1190] = 10'd9;
  assign mem[1191] = 10'd8;
  assign mem[1192] = 10'd9;
  assign mem[1193] = 10'd10;
  assign mem[1194] = 10'd11;
  assign mem[1195] = 10'd12;
  assign mem[1196] = 10'd13;
  assign mem[1197] = 10'd14;
  assign mem[1198] = 10'd15;
  assign mem[1199] = 10'd16;
  assign mem[1200] = 10'd3;
  assign mem[1201] = 10'd2;
  assign mem[1202] = 10'd1;
  assign mem[1203] = 10'd2;
  assign mem[1204] = 10'd3;
  assign mem[1205] = 10'd4;
  assign mem[1206] = 10'd5;
  assign mem[1207] = 10'd6;
  assign mem[1208] = 10'd7;
  assign mem[1209] = 10'd8;
  assign mem[1210] = 10'd2;
  assign mem[1211] = 10'd1;
  assign mem[1212] = 10'd0;
  assign mem[1213] = 10'd1;
  assign mem[1214] = 10'd2;
  assign mem[1215] = 10'd3;
  assign mem[1216] = 10'd4;
  assign mem[1217] = 10'd5;
  assign mem[1218] = 10'd6;
  assign mem[1219] = 10'd7;
  assign mem[1220] = 10'd3;
  assign mem[1221] = 10'd2;
  assign mem[1222] = 10'd1;
  assign mem[1223] = 10'd2;
  assign mem[1224] = 10'd3;
  assign mem[1225] = 10'd4;
  assign mem[1226] = 10'd5;
  assign mem[1227] = 10'd6;
  assign mem[1228] = 10'd7;
  assign mem[1229] = 10'd8;
  assign mem[1230] = 10'd4;
  assign mem[1231] = 10'd3;
  assign mem[1232] = 10'd2;
  assign mem[1233] = 10'd3;
  assign mem[1234] = 10'd4;
  assign mem[1235] = 10'd5;
  assign mem[1236] = 10'd6;
  assign mem[1237] = 10'd7;
  assign mem[1238] = 10'd8;
  assign mem[1239] = 10'd9;
  assign mem[1240] = 10'd5;
  assign mem[1241] = 10'd4;
  assign mem[1242] = 10'd3;
  assign mem[1243] = 10'd4;
  assign mem[1244] = 10'd5;
  assign mem[1245] = 10'd6;
  assign mem[1246] = 10'd7;
  assign mem[1247] = 10'd8;
  assign mem[1248] = 10'd9;
  assign mem[1249] = 10'd10;
  assign mem[1250] = 10'd6;
  assign mem[1251] = 10'd5;
  assign mem[1252] = 10'd4;
  assign mem[1253] = 10'd5;
  assign mem[1254] = 10'd6;
  assign mem[1255] = 10'd7;
  assign mem[1256] = 10'd8;
  assign mem[1257] = 10'd9;
  assign mem[1258] = 10'd10;
  assign mem[1259] = 10'd11;
  assign mem[1260] = 10'd7;
  assign mem[1261] = 10'd6;
  assign mem[1262] = 10'd5;
  assign mem[1263] = 10'd6;
  assign mem[1264] = 10'd7;
  assign mem[1265] = 10'd8;
  assign mem[1266] = 10'd9;
  assign mem[1267] = 10'd10;
  assign mem[1268] = 10'd11;
  assign mem[1269] = 10'd12;
  assign mem[1270] = 10'd8;
  assign mem[1271] = 10'd7;
  assign mem[1272] = 10'd6;
  assign mem[1273] = 10'd7;
  assign mem[1274] = 10'd8;
  assign mem[1275] = 10'd9;
  assign mem[1276] = 10'd10;
  assign mem[1277] = 10'd11;
  assign mem[1278] = 10'd12;
  assign mem[1279] = 10'd13;
  assign mem[1280] = 10'd9;
  assign mem[1281] = 10'd8;
  assign mem[1282] = 10'd7;
  assign mem[1283] = 10'd8;
  assign mem[1284] = 10'd9;
  assign mem[1285] = 10'd10;
  assign mem[1286] = 10'd11;
  assign mem[1287] = 10'd12;
  assign mem[1288] = 10'd13;
  assign mem[1289] = 10'd14;
  assign mem[1290] = 10'd10;
  assign mem[1291] = 10'd9;
  assign mem[1292] = 10'd8;
  assign mem[1293] = 10'd9;
  assign mem[1294] = 10'd10;
  assign mem[1295] = 10'd11;
  assign mem[1296] = 10'd12;
  assign mem[1297] = 10'd13;
  assign mem[1298] = 10'd14;
  assign mem[1299] = 10'd15;
  assign mem[1300] = 10'd4;
  assign mem[1301] = 10'd3;
  assign mem[1302] = 10'd2;
  assign mem[1303] = 10'd1;
  assign mem[1304] = 10'd2;
  assign mem[1305] = 10'd3;
  assign mem[1306] = 10'd4;
  assign mem[1307] = 10'd5;
  assign mem[1308] = 10'd6;
  assign mem[1309] = 10'd7;
  assign mem[1310] = 10'd3;
  assign mem[1311] = 10'd2;
  assign mem[1312] = 10'd1;
  assign mem[1313] = 10'd0;
  assign mem[1314] = 10'd1;
  assign mem[1315] = 10'd2;
  assign mem[1316] = 10'd3;
  assign mem[1317] = 10'd4;
  assign mem[1318] = 10'd5;
  assign mem[1319] = 10'd6;
  assign mem[1320] = 10'd4;
  assign mem[1321] = 10'd3;
  assign mem[1322] = 10'd2;
  assign mem[1323] = 10'd1;
  assign mem[1324] = 10'd2;
  assign mem[1325] = 10'd3;
  assign mem[1326] = 10'd4;
  assign mem[1327] = 10'd5;
  assign mem[1328] = 10'd6;
  assign mem[1329] = 10'd7;
  assign mem[1330] = 10'd5;
  assign mem[1331] = 10'd4;
  assign mem[1332] = 10'd3;
  assign mem[1333] = 10'd2;
  assign mem[1334] = 10'd3;
  assign mem[1335] = 10'd4;
  assign mem[1336] = 10'd5;
  assign mem[1337] = 10'd6;
  assign mem[1338] = 10'd7;
  assign mem[1339] = 10'd8;
  assign mem[1340] = 10'd6;
  assign mem[1341] = 10'd5;
  assign mem[1342] = 10'd4;
  assign mem[1343] = 10'd3;
  assign mem[1344] = 10'd4;
  assign mem[1345] = 10'd5;
  assign mem[1346] = 10'd6;
  assign mem[1347] = 10'd7;
  assign mem[1348] = 10'd8;
  assign mem[1349] = 10'd9;
  assign mem[1350] = 10'd7;
  assign mem[1351] = 10'd6;
  assign mem[1352] = 10'd5;
  assign mem[1353] = 10'd4;
  assign mem[1354] = 10'd5;
  assign mem[1355] = 10'd6;
  assign mem[1356] = 10'd7;
  assign mem[1357] = 10'd8;
  assign mem[1358] = 10'd9;
  assign mem[1359] = 10'd10;
  assign mem[1360] = 10'd8;
  assign mem[1361] = 10'd7;
  assign mem[1362] = 10'd6;
  assign mem[1363] = 10'd5;
  assign mem[1364] = 10'd6;
  assign mem[1365] = 10'd7;
  assign mem[1366] = 10'd8;
  assign mem[1367] = 10'd9;
  assign mem[1368] = 10'd10;
  assign mem[1369] = 10'd11;
  assign mem[1370] = 10'd9;
  assign mem[1371] = 10'd8;
  assign mem[1372] = 10'd7;
  assign mem[1373] = 10'd6;
  assign mem[1374] = 10'd7;
  assign mem[1375] = 10'd8;
  assign mem[1376] = 10'd9;
  assign mem[1377] = 10'd10;
  assign mem[1378] = 10'd11;
  assign mem[1379] = 10'd12;
  assign mem[1380] = 10'd10;
  assign mem[1381] = 10'd9;
  assign mem[1382] = 10'd8;
  assign mem[1383] = 10'd7;
  assign mem[1384] = 10'd8;
  assign mem[1385] = 10'd9;
  assign mem[1386] = 10'd10;
  assign mem[1387] = 10'd11;
  assign mem[1388] = 10'd12;
  assign mem[1389] = 10'd13;
  assign mem[1390] = 10'd11;
  assign mem[1391] = 10'd10;
  assign mem[1392] = 10'd9;
  assign mem[1393] = 10'd8;
  assign mem[1394] = 10'd9;
  assign mem[1395] = 10'd10;
  assign mem[1396] = 10'd11;
  assign mem[1397] = 10'd12;
  assign mem[1398] = 10'd13;
  assign mem[1399] = 10'd14;
  assign mem[1400] = 10'd5;
  assign mem[1401] = 10'd4;
  assign mem[1402] = 10'd3;
  assign mem[1403] = 10'd2;
  assign mem[1404] = 10'd1;
  assign mem[1405] = 10'd2;
  assign mem[1406] = 10'd3;
  assign mem[1407] = 10'd4;
  assign mem[1408] = 10'd5;
  assign mem[1409] = 10'd6;
  assign mem[1410] = 10'd4;
  assign mem[1411] = 10'd3;
  assign mem[1412] = 10'd2;
  assign mem[1413] = 10'd1;
  assign mem[1414] = 10'd0;
  assign mem[1415] = 10'd1;
  assign mem[1416] = 10'd2;
  assign mem[1417] = 10'd3;
  assign mem[1418] = 10'd4;
  assign mem[1419] = 10'd5;
  assign mem[1420] = 10'd5;
  assign mem[1421] = 10'd4;
  assign mem[1422] = 10'd3;
  assign mem[1423] = 10'd2;
  assign mem[1424] = 10'd1;
  assign mem[1425] = 10'd2;
  assign mem[1426] = 10'd3;
  assign mem[1427] = 10'd4;
  assign mem[1428] = 10'd5;
  assign mem[1429] = 10'd6;
  assign mem[1430] = 10'd6;
  assign mem[1431] = 10'd5;
  assign mem[1432] = 10'd4;
  assign mem[1433] = 10'd3;
  assign mem[1434] = 10'd2;
  assign mem[1435] = 10'd3;
  assign mem[1436] = 10'd4;
  assign mem[1437] = 10'd5;
  assign mem[1438] = 10'd6;
  assign mem[1439] = 10'd7;
  assign mem[1440] = 10'd7;
  assign mem[1441] = 10'd6;
  assign mem[1442] = 10'd5;
  assign mem[1443] = 10'd4;
  assign mem[1444] = 10'd3;
  assign mem[1445] = 10'd4;
  assign mem[1446] = 10'd5;
  assign mem[1447] = 10'd6;
  assign mem[1448] = 10'd7;
  assign mem[1449] = 10'd8;
  assign mem[1450] = 10'd8;
  assign mem[1451] = 10'd7;
  assign mem[1452] = 10'd6;
  assign mem[1453] = 10'd5;
  assign mem[1454] = 10'd4;
  assign mem[1455] = 10'd5;
  assign mem[1456] = 10'd6;
  assign mem[1457] = 10'd7;
  assign mem[1458] = 10'd8;
  assign mem[1459] = 10'd9;
  assign mem[1460] = 10'd9;
  assign mem[1461] = 10'd8;
  assign mem[1462] = 10'd7;
  assign mem[1463] = 10'd6;
  assign mem[1464] = 10'd5;
  assign mem[1465] = 10'd6;
  assign mem[1466] = 10'd7;
  assign mem[1467] = 10'd8;
  assign mem[1468] = 10'd9;
  assign mem[1469] = 10'd10;
  assign mem[1470] = 10'd10;
  assign mem[1471] = 10'd9;
  assign mem[1472] = 10'd8;
  assign mem[1473] = 10'd7;
  assign mem[1474] = 10'd6;
  assign mem[1475] = 10'd7;
  assign mem[1476] = 10'd8;
  assign mem[1477] = 10'd9;
  assign mem[1478] = 10'd10;
  assign mem[1479] = 10'd11;
  assign mem[1480] = 10'd11;
  assign mem[1481] = 10'd10;
  assign mem[1482] = 10'd9;
  assign mem[1483] = 10'd8;
  assign mem[1484] = 10'd7;
  assign mem[1485] = 10'd8;
  assign mem[1486] = 10'd9;
  assign mem[1487] = 10'd10;
  assign mem[1488] = 10'd11;
  assign mem[1489] = 10'd12;
  assign mem[1490] = 10'd12;
  assign mem[1491] = 10'd11;
  assign mem[1492] = 10'd10;
  assign mem[1493] = 10'd9;
  assign mem[1494] = 10'd8;
  assign mem[1495] = 10'd9;
  assign mem[1496] = 10'd10;
  assign mem[1497] = 10'd11;
  assign mem[1498] = 10'd12;
  assign mem[1499] = 10'd13;
  assign mem[1500] = 10'd6;
  assign mem[1501] = 10'd5;
  assign mem[1502] = 10'd4;
  assign mem[1503] = 10'd3;
  assign mem[1504] = 10'd2;
  assign mem[1505] = 10'd1;
  assign mem[1506] = 10'd2;
  assign mem[1507] = 10'd3;
  assign mem[1508] = 10'd4;
  assign mem[1509] = 10'd5;
  assign mem[1510] = 10'd5;
  assign mem[1511] = 10'd4;
  assign mem[1512] = 10'd3;
  assign mem[1513] = 10'd2;
  assign mem[1514] = 10'd1;
  assign mem[1515] = 10'd0;
  assign mem[1516] = 10'd1;
  assign mem[1517] = 10'd2;
  assign mem[1518] = 10'd3;
  assign mem[1519] = 10'd4;
  assign mem[1520] = 10'd6;
  assign mem[1521] = 10'd5;
  assign mem[1522] = 10'd4;
  assign mem[1523] = 10'd3;
  assign mem[1524] = 10'd2;
  assign mem[1525] = 10'd1;
  assign mem[1526] = 10'd2;
  assign mem[1527] = 10'd3;
  assign mem[1528] = 10'd4;
  assign mem[1529] = 10'd5;
  assign mem[1530] = 10'd7;
  assign mem[1531] = 10'd6;
  assign mem[1532] = 10'd5;
  assign mem[1533] = 10'd4;
  assign mem[1534] = 10'd3;
  assign mem[1535] = 10'd2;
  assign mem[1536] = 10'd3;
  assign mem[1537] = 10'd4;
  assign mem[1538] = 10'd5;
  assign mem[1539] = 10'd6;
  assign mem[1540] = 10'd8;
  assign mem[1541] = 10'd7;
  assign mem[1542] = 10'd6;
  assign mem[1543] = 10'd5;
  assign mem[1544] = 10'd4;
  assign mem[1545] = 10'd3;
  assign mem[1546] = 10'd4;
  assign mem[1547] = 10'd5;
  assign mem[1548] = 10'd6;
  assign mem[1549] = 10'd7;
  assign mem[1550] = 10'd9;
  assign mem[1551] = 10'd8;
  assign mem[1552] = 10'd7;
  assign mem[1553] = 10'd6;
  assign mem[1554] = 10'd5;
  assign mem[1555] = 10'd4;
  assign mem[1556] = 10'd5;
  assign mem[1557] = 10'd6;
  assign mem[1558] = 10'd7;
  assign mem[1559] = 10'd8;
  assign mem[1560] = 10'd10;
  assign mem[1561] = 10'd9;
  assign mem[1562] = 10'd8;
  assign mem[1563] = 10'd7;
  assign mem[1564] = 10'd6;
  assign mem[1565] = 10'd5;
  assign mem[1566] = 10'd6;
  assign mem[1567] = 10'd7;
  assign mem[1568] = 10'd8;
  assign mem[1569] = 10'd9;
  assign mem[1570] = 10'd11;
  assign mem[1571] = 10'd10;
  assign mem[1572] = 10'd9;
  assign mem[1573] = 10'd8;
  assign mem[1574] = 10'd7;
  assign mem[1575] = 10'd6;
  assign mem[1576] = 10'd7;
  assign mem[1577] = 10'd8;
  assign mem[1578] = 10'd9;
  assign mem[1579] = 10'd10;
  assign mem[1580] = 10'd12;
  assign mem[1581] = 10'd11;
  assign mem[1582] = 10'd10;
  assign mem[1583] = 10'd9;
  assign mem[1584] = 10'd8;
  assign mem[1585] = 10'd7;
  assign mem[1586] = 10'd8;
  assign mem[1587] = 10'd9;
  assign mem[1588] = 10'd10;
  assign mem[1589] = 10'd11;
  assign mem[1590] = 10'd13;
  assign mem[1591] = 10'd12;
  assign mem[1592] = 10'd11;
  assign mem[1593] = 10'd10;
  assign mem[1594] = 10'd9;
  assign mem[1595] = 10'd8;
  assign mem[1596] = 10'd9;
  assign mem[1597] = 10'd10;
  assign mem[1598] = 10'd11;
  assign mem[1599] = 10'd12;
  assign mem[1600] = 10'd7;
  assign mem[1601] = 10'd6;
  assign mem[1602] = 10'd5;
  assign mem[1603] = 10'd4;
  assign mem[1604] = 10'd3;
  assign mem[1605] = 10'd2;
  assign mem[1606] = 10'd1;
  assign mem[1607] = 10'd2;
  assign mem[1608] = 10'd3;
  assign mem[1609] = 10'd4;
  assign mem[1610] = 10'd6;
  assign mem[1611] = 10'd5;
  assign mem[1612] = 10'd4;
  assign mem[1613] = 10'd3;
  assign mem[1614] = 10'd2;
  assign mem[1615] = 10'd1;
  assign mem[1616] = 10'd0;
  assign mem[1617] = 10'd1;
  assign mem[1618] = 10'd2;
  assign mem[1619] = 10'd3;
  assign mem[1620] = 10'd7;
  assign mem[1621] = 10'd6;
  assign mem[1622] = 10'd5;
  assign mem[1623] = 10'd4;
  assign mem[1624] = 10'd3;
  assign mem[1625] = 10'd2;
  assign mem[1626] = 10'd1;
  assign mem[1627] = 10'd2;
  assign mem[1628] = 10'd3;
  assign mem[1629] = 10'd4;
  assign mem[1630] = 10'd8;
  assign mem[1631] = 10'd7;
  assign mem[1632] = 10'd6;
  assign mem[1633] = 10'd5;
  assign mem[1634] = 10'd4;
  assign mem[1635] = 10'd3;
  assign mem[1636] = 10'd2;
  assign mem[1637] = 10'd3;
  assign mem[1638] = 10'd4;
  assign mem[1639] = 10'd5;
  assign mem[1640] = 10'd9;
  assign mem[1641] = 10'd8;
  assign mem[1642] = 10'd7;
  assign mem[1643] = 10'd6;
  assign mem[1644] = 10'd5;
  assign mem[1645] = 10'd4;
  assign mem[1646] = 10'd3;
  assign mem[1647] = 10'd4;
  assign mem[1648] = 10'd5;
  assign mem[1649] = 10'd6;
  assign mem[1650] = 10'd10;
  assign mem[1651] = 10'd9;
  assign mem[1652] = 10'd8;
  assign mem[1653] = 10'd7;
  assign mem[1654] = 10'd6;
  assign mem[1655] = 10'd5;
  assign mem[1656] = 10'd4;
  assign mem[1657] = 10'd5;
  assign mem[1658] = 10'd6;
  assign mem[1659] = 10'd7;
  assign mem[1660] = 10'd11;
  assign mem[1661] = 10'd10;
  assign mem[1662] = 10'd9;
  assign mem[1663] = 10'd8;
  assign mem[1664] = 10'd7;
  assign mem[1665] = 10'd6;
  assign mem[1666] = 10'd5;
  assign mem[1667] = 10'd6;
  assign mem[1668] = 10'd7;
  assign mem[1669] = 10'd8;
  assign mem[1670] = 10'd12;
  assign mem[1671] = 10'd11;
  assign mem[1672] = 10'd10;
  assign mem[1673] = 10'd9;
  assign mem[1674] = 10'd8;
  assign mem[1675] = 10'd7;
  assign mem[1676] = 10'd6;
  assign mem[1677] = 10'd7;
  assign mem[1678] = 10'd8;
  assign mem[1679] = 10'd9;
  assign mem[1680] = 10'd13;
  assign mem[1681] = 10'd12;
  assign mem[1682] = 10'd11;
  assign mem[1683] = 10'd10;
  assign mem[1684] = 10'd9;
  assign mem[1685] = 10'd8;
  assign mem[1686] = 10'd7;
  assign mem[1687] = 10'd8;
  assign mem[1688] = 10'd9;
  assign mem[1689] = 10'd10;
  assign mem[1690] = 10'd14;
  assign mem[1691] = 10'd13;
  assign mem[1692] = 10'd12;
  assign mem[1693] = 10'd11;
  assign mem[1694] = 10'd10;
  assign mem[1695] = 10'd9;
  assign mem[1696] = 10'd8;
  assign mem[1697] = 10'd9;
  assign mem[1698] = 10'd10;
  assign mem[1699] = 10'd11;
  assign mem[1700] = 10'd8;
  assign mem[1701] = 10'd7;
  assign mem[1702] = 10'd6;
  assign mem[1703] = 10'd5;
  assign mem[1704] = 10'd4;
  assign mem[1705] = 10'd3;
  assign mem[1706] = 10'd2;
  assign mem[1707] = 10'd1;
  assign mem[1708] = 10'd2;
  assign mem[1709] = 10'd3;
  assign mem[1710] = 10'd7;
  assign mem[1711] = 10'd6;
  assign mem[1712] = 10'd5;
  assign mem[1713] = 10'd4;
  assign mem[1714] = 10'd3;
  assign mem[1715] = 10'd2;
  assign mem[1716] = 10'd1;
  assign mem[1717] = 10'd0;
  assign mem[1718] = 10'd1;
  assign mem[1719] = 10'd2;
  assign mem[1720] = 10'd8;
  assign mem[1721] = 10'd7;
  assign mem[1722] = 10'd6;
  assign mem[1723] = 10'd5;
  assign mem[1724] = 10'd4;
  assign mem[1725] = 10'd3;
  assign mem[1726] = 10'd2;
  assign mem[1727] = 10'd1;
  assign mem[1728] = 10'd2;
  assign mem[1729] = 10'd3;
  assign mem[1730] = 10'd9;
  assign mem[1731] = 10'd8;
  assign mem[1732] = 10'd7;
  assign mem[1733] = 10'd6;
  assign mem[1734] = 10'd5;
  assign mem[1735] = 10'd4;
  assign mem[1736] = 10'd3;
  assign mem[1737] = 10'd2;
  assign mem[1738] = 10'd3;
  assign mem[1739] = 10'd4;
  assign mem[1740] = 10'd10;
  assign mem[1741] = 10'd9;
  assign mem[1742] = 10'd8;
  assign mem[1743] = 10'd7;
  assign mem[1744] = 10'd6;
  assign mem[1745] = 10'd5;
  assign mem[1746] = 10'd4;
  assign mem[1747] = 10'd3;
  assign mem[1748] = 10'd4;
  assign mem[1749] = 10'd5;
  assign mem[1750] = 10'd11;
  assign mem[1751] = 10'd10;
  assign mem[1752] = 10'd9;
  assign mem[1753] = 10'd8;
  assign mem[1754] = 10'd7;
  assign mem[1755] = 10'd6;
  assign mem[1756] = 10'd5;
  assign mem[1757] = 10'd4;
  assign mem[1758] = 10'd5;
  assign mem[1759] = 10'd6;
  assign mem[1760] = 10'd12;
  assign mem[1761] = 10'd11;
  assign mem[1762] = 10'd10;
  assign mem[1763] = 10'd9;
  assign mem[1764] = 10'd8;
  assign mem[1765] = 10'd7;
  assign mem[1766] = 10'd6;
  assign mem[1767] = 10'd5;
  assign mem[1768] = 10'd6;
  assign mem[1769] = 10'd7;
  assign mem[1770] = 10'd13;
  assign mem[1771] = 10'd12;
  assign mem[1772] = 10'd11;
  assign mem[1773] = 10'd10;
  assign mem[1774] = 10'd9;
  assign mem[1775] = 10'd8;
  assign mem[1776] = 10'd7;
  assign mem[1777] = 10'd6;
  assign mem[1778] = 10'd7;
  assign mem[1779] = 10'd8;
  assign mem[1780] = 10'd14;
  assign mem[1781] = 10'd13;
  assign mem[1782] = 10'd12;
  assign mem[1783] = 10'd11;
  assign mem[1784] = 10'd10;
  assign mem[1785] = 10'd9;
  assign mem[1786] = 10'd8;
  assign mem[1787] = 10'd7;
  assign mem[1788] = 10'd8;
  assign mem[1789] = 10'd9;
  assign mem[1790] = 10'd15;
  assign mem[1791] = 10'd14;
  assign mem[1792] = 10'd13;
  assign mem[1793] = 10'd12;
  assign mem[1794] = 10'd11;
  assign mem[1795] = 10'd10;
  assign mem[1796] = 10'd9;
  assign mem[1797] = 10'd8;
  assign mem[1798] = 10'd9;
  assign mem[1799] = 10'd10;
  assign mem[1800] = 10'd9;
  assign mem[1801] = 10'd8;
  assign mem[1802] = 10'd7;
  assign mem[1803] = 10'd6;
  assign mem[1804] = 10'd5;
  assign mem[1805] = 10'd4;
  assign mem[1806] = 10'd3;
  assign mem[1807] = 10'd2;
  assign mem[1808] = 10'd1;
  assign mem[1809] = 10'd2;
  assign mem[1810] = 10'd8;
  assign mem[1811] = 10'd7;
  assign mem[1812] = 10'd6;
  assign mem[1813] = 10'd5;
  assign mem[1814] = 10'd4;
  assign mem[1815] = 10'd3;
  assign mem[1816] = 10'd2;
  assign mem[1817] = 10'd1;
  assign mem[1818] = 10'd0;
  assign mem[1819] = 10'd1;
  assign mem[1820] = 10'd9;
  assign mem[1821] = 10'd8;
  assign mem[1822] = 10'd7;
  assign mem[1823] = 10'd6;
  assign mem[1824] = 10'd5;
  assign mem[1825] = 10'd4;
  assign mem[1826] = 10'd3;
  assign mem[1827] = 10'd2;
  assign mem[1828] = 10'd1;
  assign mem[1829] = 10'd2;
  assign mem[1830] = 10'd10;
  assign mem[1831] = 10'd9;
  assign mem[1832] = 10'd8;
  assign mem[1833] = 10'd7;
  assign mem[1834] = 10'd6;
  assign mem[1835] = 10'd5;
  assign mem[1836] = 10'd4;
  assign mem[1837] = 10'd3;
  assign mem[1838] = 10'd2;
  assign mem[1839] = 10'd3;
  assign mem[1840] = 10'd11;
  assign mem[1841] = 10'd10;
  assign mem[1842] = 10'd9;
  assign mem[1843] = 10'd8;
  assign mem[1844] = 10'd7;
  assign mem[1845] = 10'd6;
  assign mem[1846] = 10'd5;
  assign mem[1847] = 10'd4;
  assign mem[1848] = 10'd3;
  assign mem[1849] = 10'd4;
  assign mem[1850] = 10'd12;
  assign mem[1851] = 10'd11;
  assign mem[1852] = 10'd10;
  assign mem[1853] = 10'd9;
  assign mem[1854] = 10'd8;
  assign mem[1855] = 10'd7;
  assign mem[1856] = 10'd6;
  assign mem[1857] = 10'd5;
  assign mem[1858] = 10'd4;
  assign mem[1859] = 10'd5;
  assign mem[1860] = 10'd13;
  assign mem[1861] = 10'd12;
  assign mem[1862] = 10'd11;
  assign mem[1863] = 10'd10;
  assign mem[1864] = 10'd9;
  assign mem[1865] = 10'd8;
  assign mem[1866] = 10'd7;
  assign mem[1867] = 10'd6;
  assign mem[1868] = 10'd5;
  assign mem[1869] = 10'd6;
  assign mem[1870] = 10'd14;
  assign mem[1871] = 10'd13;
  assign mem[1872] = 10'd12;
  assign mem[1873] = 10'd11;
  assign mem[1874] = 10'd10;
  assign mem[1875] = 10'd9;
  assign mem[1876] = 10'd8;
  assign mem[1877] = 10'd7;
  assign mem[1878] = 10'd6;
  assign mem[1879] = 10'd7;
  assign mem[1880] = 10'd15;
  assign mem[1881] = 10'd14;
  assign mem[1882] = 10'd13;
  assign mem[1883] = 10'd12;
  assign mem[1884] = 10'd11;
  assign mem[1885] = 10'd10;
  assign mem[1886] = 10'd9;
  assign mem[1887] = 10'd8;
  assign mem[1888] = 10'd7;
  assign mem[1889] = 10'd8;
  assign mem[1890] = 10'd16;
  assign mem[1891] = 10'd15;
  assign mem[1892] = 10'd14;
  assign mem[1893] = 10'd13;
  assign mem[1894] = 10'd12;
  assign mem[1895] = 10'd11;
  assign mem[1896] = 10'd10;
  assign mem[1897] = 10'd9;
  assign mem[1898] = 10'd8;
  assign mem[1899] = 10'd9;
  assign mem[1900] = 10'd10;
  assign mem[1901] = 10'd9;
  assign mem[1902] = 10'd8;
  assign mem[1903] = 10'd7;
  assign mem[1904] = 10'd6;
  assign mem[1905] = 10'd5;
  assign mem[1906] = 10'd4;
  assign mem[1907] = 10'd3;
  assign mem[1908] = 10'd2;
  assign mem[1909] = 10'd1;
  assign mem[1910] = 10'd9;
  assign mem[1911] = 10'd8;
  assign mem[1912] = 10'd7;
  assign mem[1913] = 10'd6;
  assign mem[1914] = 10'd5;
  assign mem[1915] = 10'd4;
  assign mem[1916] = 10'd3;
  assign mem[1917] = 10'd2;
  assign mem[1918] = 10'd1;
  assign mem[1919] = 10'd0;
  assign mem[1920] = 10'd10;
  assign mem[1921] = 10'd9;
  assign mem[1922] = 10'd8;
  assign mem[1923] = 10'd7;
  assign mem[1924] = 10'd6;
  assign mem[1925] = 10'd5;
  assign mem[1926] = 10'd4;
  assign mem[1927] = 10'd3;
  assign mem[1928] = 10'd2;
  assign mem[1929] = 10'd1;
  assign mem[1930] = 10'd11;
  assign mem[1931] = 10'd10;
  assign mem[1932] = 10'd9;
  assign mem[1933] = 10'd8;
  assign mem[1934] = 10'd7;
  assign mem[1935] = 10'd6;
  assign mem[1936] = 10'd5;
  assign mem[1937] = 10'd4;
  assign mem[1938] = 10'd3;
  assign mem[1939] = 10'd2;
  assign mem[1940] = 10'd12;
  assign mem[1941] = 10'd11;
  assign mem[1942] = 10'd10;
  assign mem[1943] = 10'd9;
  assign mem[1944] = 10'd8;
  assign mem[1945] = 10'd7;
  assign mem[1946] = 10'd6;
  assign mem[1947] = 10'd5;
  assign mem[1948] = 10'd4;
  assign mem[1949] = 10'd3;
  assign mem[1950] = 10'd13;
  assign mem[1951] = 10'd12;
  assign mem[1952] = 10'd11;
  assign mem[1953] = 10'd10;
  assign mem[1954] = 10'd9;
  assign mem[1955] = 10'd8;
  assign mem[1956] = 10'd7;
  assign mem[1957] = 10'd6;
  assign mem[1958] = 10'd5;
  assign mem[1959] = 10'd4;
  assign mem[1960] = 10'd14;
  assign mem[1961] = 10'd13;
  assign mem[1962] = 10'd12;
  assign mem[1963] = 10'd11;
  assign mem[1964] = 10'd10;
  assign mem[1965] = 10'd9;
  assign mem[1966] = 10'd8;
  assign mem[1967] = 10'd7;
  assign mem[1968] = 10'd6;
  assign mem[1969] = 10'd5;
  assign mem[1970] = 10'd15;
  assign mem[1971] = 10'd14;
  assign mem[1972] = 10'd13;
  assign mem[1973] = 10'd12;
  assign mem[1974] = 10'd11;
  assign mem[1975] = 10'd10;
  assign mem[1976] = 10'd9;
  assign mem[1977] = 10'd8;
  assign mem[1978] = 10'd7;
  assign mem[1979] = 10'd6;
  assign mem[1980] = 10'd16;
  assign mem[1981] = 10'd15;
  assign mem[1982] = 10'd14;
  assign mem[1983] = 10'd13;
  assign mem[1984] = 10'd12;
  assign mem[1985] = 10'd11;
  assign mem[1986] = 10'd10;
  assign mem[1987] = 10'd9;
  assign mem[1988] = 10'd8;
  assign mem[1989] = 10'd7;
  assign mem[1990] = 10'd17;
  assign mem[1991] = 10'd16;
  assign mem[1992] = 10'd15;
  assign mem[1993] = 10'd14;
  assign mem[1994] = 10'd13;
  assign mem[1995] = 10'd12;
  assign mem[1996] = 10'd11;
  assign mem[1997] = 10'd10;
  assign mem[1998] = 10'd9;
  assign mem[1999] = 10'd8;
  assign mem[2000] = 10'd2;
  assign mem[2001] = 10'd3;
  assign mem[2002] = 10'd4;
  assign mem[2003] = 10'd5;
  assign mem[2004] = 10'd6;
  assign mem[2005] = 10'd7;
  assign mem[2006] = 10'd8;
  assign mem[2007] = 10'd9;
  assign mem[2008] = 10'd10;
  assign mem[2009] = 10'd11;
  assign mem[2010] = 10'd1;
  assign mem[2011] = 10'd2;
  assign mem[2012] = 10'd3;
  assign mem[2013] = 10'd4;
  assign mem[2014] = 10'd5;
  assign mem[2015] = 10'd6;
  assign mem[2016] = 10'd7;
  assign mem[2017] = 10'd8;
  assign mem[2018] = 10'd9;
  assign mem[2019] = 10'd10;
  assign mem[2020] = 10'd0;
  assign mem[2021] = 10'd1;
  assign mem[2022] = 10'd2;
  assign mem[2023] = 10'd3;
  assign mem[2024] = 10'd4;
  assign mem[2025] = 10'd5;
  assign mem[2026] = 10'd6;
  assign mem[2027] = 10'd7;
  assign mem[2028] = 10'd8;
  assign mem[2029] = 10'd9;
  assign mem[2030] = 10'd1;
  assign mem[2031] = 10'd2;
  assign mem[2032] = 10'd3;
  assign mem[2033] = 10'd4;
  assign mem[2034] = 10'd5;
  assign mem[2035] = 10'd6;
  assign mem[2036] = 10'd7;
  assign mem[2037] = 10'd8;
  assign mem[2038] = 10'd9;
  assign mem[2039] = 10'd10;
  assign mem[2040] = 10'd2;
  assign mem[2041] = 10'd3;
  assign mem[2042] = 10'd4;
  assign mem[2043] = 10'd5;
  assign mem[2044] = 10'd6;
  assign mem[2045] = 10'd7;
  assign mem[2046] = 10'd8;
  assign mem[2047] = 10'd9;
  assign mem[2048] = 10'd10;
  assign mem[2049] = 10'd11;
  assign mem[2050] = 10'd3;
  assign mem[2051] = 10'd4;
  assign mem[2052] = 10'd5;
  assign mem[2053] = 10'd6;
  assign mem[2054] = 10'd7;
  assign mem[2055] = 10'd8;
  assign mem[2056] = 10'd9;
  assign mem[2057] = 10'd10;
  assign mem[2058] = 10'd11;
  assign mem[2059] = 10'd12;
  assign mem[2060] = 10'd4;
  assign mem[2061] = 10'd5;
  assign mem[2062] = 10'd6;
  assign mem[2063] = 10'd7;
  assign mem[2064] = 10'd8;
  assign mem[2065] = 10'd9;
  assign mem[2066] = 10'd10;
  assign mem[2067] = 10'd11;
  assign mem[2068] = 10'd12;
  assign mem[2069] = 10'd13;
  assign mem[2070] = 10'd5;
  assign mem[2071] = 10'd6;
  assign mem[2072] = 10'd7;
  assign mem[2073] = 10'd8;
  assign mem[2074] = 10'd9;
  assign mem[2075] = 10'd10;
  assign mem[2076] = 10'd11;
  assign mem[2077] = 10'd12;
  assign mem[2078] = 10'd13;
  assign mem[2079] = 10'd14;
  assign mem[2080] = 10'd6;
  assign mem[2081] = 10'd7;
  assign mem[2082] = 10'd8;
  assign mem[2083] = 10'd9;
  assign mem[2084] = 10'd10;
  assign mem[2085] = 10'd11;
  assign mem[2086] = 10'd12;
  assign mem[2087] = 10'd13;
  assign mem[2088] = 10'd14;
  assign mem[2089] = 10'd15;
  assign mem[2090] = 10'd7;
  assign mem[2091] = 10'd8;
  assign mem[2092] = 10'd9;
  assign mem[2093] = 10'd10;
  assign mem[2094] = 10'd11;
  assign mem[2095] = 10'd12;
  assign mem[2096] = 10'd13;
  assign mem[2097] = 10'd14;
  assign mem[2098] = 10'd15;
  assign mem[2099] = 10'd16;
  assign mem[2100] = 10'd3;
  assign mem[2101] = 10'd2;
  assign mem[2102] = 10'd3;
  assign mem[2103] = 10'd4;
  assign mem[2104] = 10'd5;
  assign mem[2105] = 10'd6;
  assign mem[2106] = 10'd7;
  assign mem[2107] = 10'd8;
  assign mem[2108] = 10'd9;
  assign mem[2109] = 10'd10;
  assign mem[2110] = 10'd2;
  assign mem[2111] = 10'd1;
  assign mem[2112] = 10'd2;
  assign mem[2113] = 10'd3;
  assign mem[2114] = 10'd4;
  assign mem[2115] = 10'd5;
  assign mem[2116] = 10'd6;
  assign mem[2117] = 10'd7;
  assign mem[2118] = 10'd8;
  assign mem[2119] = 10'd9;
  assign mem[2120] = 10'd1;
  assign mem[2121] = 10'd0;
  assign mem[2122] = 10'd1;
  assign mem[2123] = 10'd2;
  assign mem[2124] = 10'd3;
  assign mem[2125] = 10'd4;
  assign mem[2126] = 10'd5;
  assign mem[2127] = 10'd6;
  assign mem[2128] = 10'd7;
  assign mem[2129] = 10'd8;
  assign mem[2130] = 10'd2;
  assign mem[2131] = 10'd1;
  assign mem[2132] = 10'd2;
  assign mem[2133] = 10'd3;
  assign mem[2134] = 10'd4;
  assign mem[2135] = 10'd5;
  assign mem[2136] = 10'd6;
  assign mem[2137] = 10'd7;
  assign mem[2138] = 10'd8;
  assign mem[2139] = 10'd9;
  assign mem[2140] = 10'd3;
  assign mem[2141] = 10'd2;
  assign mem[2142] = 10'd3;
  assign mem[2143] = 10'd4;
  assign mem[2144] = 10'd5;
  assign mem[2145] = 10'd6;
  assign mem[2146] = 10'd7;
  assign mem[2147] = 10'd8;
  assign mem[2148] = 10'd9;
  assign mem[2149] = 10'd10;
  assign mem[2150] = 10'd4;
  assign mem[2151] = 10'd3;
  assign mem[2152] = 10'd4;
  assign mem[2153] = 10'd5;
  assign mem[2154] = 10'd6;
  assign mem[2155] = 10'd7;
  assign mem[2156] = 10'd8;
  assign mem[2157] = 10'd9;
  assign mem[2158] = 10'd10;
  assign mem[2159] = 10'd11;
  assign mem[2160] = 10'd5;
  assign mem[2161] = 10'd4;
  assign mem[2162] = 10'd5;
  assign mem[2163] = 10'd6;
  assign mem[2164] = 10'd7;
  assign mem[2165] = 10'd8;
  assign mem[2166] = 10'd9;
  assign mem[2167] = 10'd10;
  assign mem[2168] = 10'd11;
  assign mem[2169] = 10'd12;
  assign mem[2170] = 10'd6;
  assign mem[2171] = 10'd5;
  assign mem[2172] = 10'd6;
  assign mem[2173] = 10'd7;
  assign mem[2174] = 10'd8;
  assign mem[2175] = 10'd9;
  assign mem[2176] = 10'd10;
  assign mem[2177] = 10'd11;
  assign mem[2178] = 10'd12;
  assign mem[2179] = 10'd13;
  assign mem[2180] = 10'd7;
  assign mem[2181] = 10'd6;
  assign mem[2182] = 10'd7;
  assign mem[2183] = 10'd8;
  assign mem[2184] = 10'd9;
  assign mem[2185] = 10'd10;
  assign mem[2186] = 10'd11;
  assign mem[2187] = 10'd12;
  assign mem[2188] = 10'd13;
  assign mem[2189] = 10'd14;
  assign mem[2190] = 10'd8;
  assign mem[2191] = 10'd7;
  assign mem[2192] = 10'd8;
  assign mem[2193] = 10'd9;
  assign mem[2194] = 10'd10;
  assign mem[2195] = 10'd11;
  assign mem[2196] = 10'd12;
  assign mem[2197] = 10'd13;
  assign mem[2198] = 10'd14;
  assign mem[2199] = 10'd15;
  assign mem[2200] = 10'd4;
  assign mem[2201] = 10'd3;
  assign mem[2202] = 10'd2;
  assign mem[2203] = 10'd3;
  assign mem[2204] = 10'd4;
  assign mem[2205] = 10'd5;
  assign mem[2206] = 10'd6;
  assign mem[2207] = 10'd7;
  assign mem[2208] = 10'd8;
  assign mem[2209] = 10'd9;
  assign mem[2210] = 10'd3;
  assign mem[2211] = 10'd2;
  assign mem[2212] = 10'd1;
  assign mem[2213] = 10'd2;
  assign mem[2214] = 10'd3;
  assign mem[2215] = 10'd4;
  assign mem[2216] = 10'd5;
  assign mem[2217] = 10'd6;
  assign mem[2218] = 10'd7;
  assign mem[2219] = 10'd8;
  assign mem[2220] = 10'd2;
  assign mem[2221] = 10'd1;
  assign mem[2222] = 10'd0;
  assign mem[2223] = 10'd1;
  assign mem[2224] = 10'd2;
  assign mem[2225] = 10'd3;
  assign mem[2226] = 10'd4;
  assign mem[2227] = 10'd5;
  assign mem[2228] = 10'd6;
  assign mem[2229] = 10'd7;
  assign mem[2230] = 10'd3;
  assign mem[2231] = 10'd2;
  assign mem[2232] = 10'd1;
  assign mem[2233] = 10'd2;
  assign mem[2234] = 10'd3;
  assign mem[2235] = 10'd4;
  assign mem[2236] = 10'd5;
  assign mem[2237] = 10'd6;
  assign mem[2238] = 10'd7;
  assign mem[2239] = 10'd8;
  assign mem[2240] = 10'd4;
  assign mem[2241] = 10'd3;
  assign mem[2242] = 10'd2;
  assign mem[2243] = 10'd3;
  assign mem[2244] = 10'd4;
  assign mem[2245] = 10'd5;
  assign mem[2246] = 10'd6;
  assign mem[2247] = 10'd7;
  assign mem[2248] = 10'd8;
  assign mem[2249] = 10'd9;
  assign mem[2250] = 10'd5;
  assign mem[2251] = 10'd4;
  assign mem[2252] = 10'd3;
  assign mem[2253] = 10'd4;
  assign mem[2254] = 10'd5;
  assign mem[2255] = 10'd6;
  assign mem[2256] = 10'd7;
  assign mem[2257] = 10'd8;
  assign mem[2258] = 10'd9;
  assign mem[2259] = 10'd10;
  assign mem[2260] = 10'd6;
  assign mem[2261] = 10'd5;
  assign mem[2262] = 10'd4;
  assign mem[2263] = 10'd5;
  assign mem[2264] = 10'd6;
  assign mem[2265] = 10'd7;
  assign mem[2266] = 10'd8;
  assign mem[2267] = 10'd9;
  assign mem[2268] = 10'd10;
  assign mem[2269] = 10'd11;
  assign mem[2270] = 10'd7;
  assign mem[2271] = 10'd6;
  assign mem[2272] = 10'd5;
  assign mem[2273] = 10'd6;
  assign mem[2274] = 10'd7;
  assign mem[2275] = 10'd8;
  assign mem[2276] = 10'd9;
  assign mem[2277] = 10'd10;
  assign mem[2278] = 10'd11;
  assign mem[2279] = 10'd12;
  assign mem[2280] = 10'd8;
  assign mem[2281] = 10'd7;
  assign mem[2282] = 10'd6;
  assign mem[2283] = 10'd7;
  assign mem[2284] = 10'd8;
  assign mem[2285] = 10'd9;
  assign mem[2286] = 10'd10;
  assign mem[2287] = 10'd11;
  assign mem[2288] = 10'd12;
  assign mem[2289] = 10'd13;
  assign mem[2290] = 10'd9;
  assign mem[2291] = 10'd8;
  assign mem[2292] = 10'd7;
  assign mem[2293] = 10'd8;
  assign mem[2294] = 10'd9;
  assign mem[2295] = 10'd10;
  assign mem[2296] = 10'd11;
  assign mem[2297] = 10'd12;
  assign mem[2298] = 10'd13;
  assign mem[2299] = 10'd14;
  assign mem[2300] = 10'd5;
  assign mem[2301] = 10'd4;
  assign mem[2302] = 10'd3;
  assign mem[2303] = 10'd2;
  assign mem[2304] = 10'd3;
  assign mem[2305] = 10'd4;
  assign mem[2306] = 10'd5;
  assign mem[2307] = 10'd6;
  assign mem[2308] = 10'd7;
  assign mem[2309] = 10'd8;
  assign mem[2310] = 10'd4;
  assign mem[2311] = 10'd3;
  assign mem[2312] = 10'd2;
  assign mem[2313] = 10'd1;
  assign mem[2314] = 10'd2;
  assign mem[2315] = 10'd3;
  assign mem[2316] = 10'd4;
  assign mem[2317] = 10'd5;
  assign mem[2318] = 10'd6;
  assign mem[2319] = 10'd7;
  assign mem[2320] = 10'd3;
  assign mem[2321] = 10'd2;
  assign mem[2322] = 10'd1;
  assign mem[2323] = 10'd0;
  assign mem[2324] = 10'd1;
  assign mem[2325] = 10'd2;
  assign mem[2326] = 10'd3;
  assign mem[2327] = 10'd4;
  assign mem[2328] = 10'd5;
  assign mem[2329] = 10'd6;
  assign mem[2330] = 10'd4;
  assign mem[2331] = 10'd3;
  assign mem[2332] = 10'd2;
  assign mem[2333] = 10'd1;
  assign mem[2334] = 10'd2;
  assign mem[2335] = 10'd3;
  assign mem[2336] = 10'd4;
  assign mem[2337] = 10'd5;
  assign mem[2338] = 10'd6;
  assign mem[2339] = 10'd7;
  assign mem[2340] = 10'd5;
  assign mem[2341] = 10'd4;
  assign mem[2342] = 10'd3;
  assign mem[2343] = 10'd2;
  assign mem[2344] = 10'd3;
  assign mem[2345] = 10'd4;
  assign mem[2346] = 10'd5;
  assign mem[2347] = 10'd6;
  assign mem[2348] = 10'd7;
  assign mem[2349] = 10'd8;
  assign mem[2350] = 10'd6;
  assign mem[2351] = 10'd5;
  assign mem[2352] = 10'd4;
  assign mem[2353] = 10'd3;
  assign mem[2354] = 10'd4;
  assign mem[2355] = 10'd5;
  assign mem[2356] = 10'd6;
  assign mem[2357] = 10'd7;
  assign mem[2358] = 10'd8;
  assign mem[2359] = 10'd9;
  assign mem[2360] = 10'd7;
  assign mem[2361] = 10'd6;
  assign mem[2362] = 10'd5;
  assign mem[2363] = 10'd4;
  assign mem[2364] = 10'd5;
  assign mem[2365] = 10'd6;
  assign mem[2366] = 10'd7;
  assign mem[2367] = 10'd8;
  assign mem[2368] = 10'd9;
  assign mem[2369] = 10'd10;
  assign mem[2370] = 10'd8;
  assign mem[2371] = 10'd7;
  assign mem[2372] = 10'd6;
  assign mem[2373] = 10'd5;
  assign mem[2374] = 10'd6;
  assign mem[2375] = 10'd7;
  assign mem[2376] = 10'd8;
  assign mem[2377] = 10'd9;
  assign mem[2378] = 10'd10;
  assign mem[2379] = 10'd11;
  assign mem[2380] = 10'd9;
  assign mem[2381] = 10'd8;
  assign mem[2382] = 10'd7;
  assign mem[2383] = 10'd6;
  assign mem[2384] = 10'd7;
  assign mem[2385] = 10'd8;
  assign mem[2386] = 10'd9;
  assign mem[2387] = 10'd10;
  assign mem[2388] = 10'd11;
  assign mem[2389] = 10'd12;
  assign mem[2390] = 10'd10;
  assign mem[2391] = 10'd9;
  assign mem[2392] = 10'd8;
  assign mem[2393] = 10'd7;
  assign mem[2394] = 10'd8;
  assign mem[2395] = 10'd9;
  assign mem[2396] = 10'd10;
  assign mem[2397] = 10'd11;
  assign mem[2398] = 10'd12;
  assign mem[2399] = 10'd13;
  assign mem[2400] = 10'd6;
  assign mem[2401] = 10'd5;
  assign mem[2402] = 10'd4;
  assign mem[2403] = 10'd3;
  assign mem[2404] = 10'd2;
  assign mem[2405] = 10'd3;
  assign mem[2406] = 10'd4;
  assign mem[2407] = 10'd5;
  assign mem[2408] = 10'd6;
  assign mem[2409] = 10'd7;
  assign mem[2410] = 10'd5;
  assign mem[2411] = 10'd4;
  assign mem[2412] = 10'd3;
  assign mem[2413] = 10'd2;
  assign mem[2414] = 10'd1;
  assign mem[2415] = 10'd2;
  assign mem[2416] = 10'd3;
  assign mem[2417] = 10'd4;
  assign mem[2418] = 10'd5;
  assign mem[2419] = 10'd6;
  assign mem[2420] = 10'd4;
  assign mem[2421] = 10'd3;
  assign mem[2422] = 10'd2;
  assign mem[2423] = 10'd1;
  assign mem[2424] = 10'd0;
  assign mem[2425] = 10'd1;
  assign mem[2426] = 10'd2;
  assign mem[2427] = 10'd3;
  assign mem[2428] = 10'd4;
  assign mem[2429] = 10'd5;
  assign mem[2430] = 10'd5;
  assign mem[2431] = 10'd4;
  assign mem[2432] = 10'd3;
  assign mem[2433] = 10'd2;
  assign mem[2434] = 10'd1;
  assign mem[2435] = 10'd2;
  assign mem[2436] = 10'd3;
  assign mem[2437] = 10'd4;
  assign mem[2438] = 10'd5;
  assign mem[2439] = 10'd6;
  assign mem[2440] = 10'd6;
  assign mem[2441] = 10'd5;
  assign mem[2442] = 10'd4;
  assign mem[2443] = 10'd3;
  assign mem[2444] = 10'd2;
  assign mem[2445] = 10'd3;
  assign mem[2446] = 10'd4;
  assign mem[2447] = 10'd5;
  assign mem[2448] = 10'd6;
  assign mem[2449] = 10'd7;
  assign mem[2450] = 10'd7;
  assign mem[2451] = 10'd6;
  assign mem[2452] = 10'd5;
  assign mem[2453] = 10'd4;
  assign mem[2454] = 10'd3;
  assign mem[2455] = 10'd4;
  assign mem[2456] = 10'd5;
  assign mem[2457] = 10'd6;
  assign mem[2458] = 10'd7;
  assign mem[2459] = 10'd8;
  assign mem[2460] = 10'd8;
  assign mem[2461] = 10'd7;
  assign mem[2462] = 10'd6;
  assign mem[2463] = 10'd5;
  assign mem[2464] = 10'd4;
  assign mem[2465] = 10'd5;
  assign mem[2466] = 10'd6;
  assign mem[2467] = 10'd7;
  assign mem[2468] = 10'd8;
  assign mem[2469] = 10'd9;
  assign mem[2470] = 10'd9;
  assign mem[2471] = 10'd8;
  assign mem[2472] = 10'd7;
  assign mem[2473] = 10'd6;
  assign mem[2474] = 10'd5;
  assign mem[2475] = 10'd6;
  assign mem[2476] = 10'd7;
  assign mem[2477] = 10'd8;
  assign mem[2478] = 10'd9;
  assign mem[2479] = 10'd10;
  assign mem[2480] = 10'd10;
  assign mem[2481] = 10'd9;
  assign mem[2482] = 10'd8;
  assign mem[2483] = 10'd7;
  assign mem[2484] = 10'd6;
  assign mem[2485] = 10'd7;
  assign mem[2486] = 10'd8;
  assign mem[2487] = 10'd9;
  assign mem[2488] = 10'd10;
  assign mem[2489] = 10'd11;
  assign mem[2490] = 10'd11;
  assign mem[2491] = 10'd10;
  assign mem[2492] = 10'd9;
  assign mem[2493] = 10'd8;
  assign mem[2494] = 10'd7;
  assign mem[2495] = 10'd8;
  assign mem[2496] = 10'd9;
  assign mem[2497] = 10'd10;
  assign mem[2498] = 10'd11;
  assign mem[2499] = 10'd12;
  assign mem[2500] = 10'd7;
  assign mem[2501] = 10'd6;
  assign mem[2502] = 10'd5;
  assign mem[2503] = 10'd4;
  assign mem[2504] = 10'd3;
  assign mem[2505] = 10'd2;
  assign mem[2506] = 10'd3;
  assign mem[2507] = 10'd4;
  assign mem[2508] = 10'd5;
  assign mem[2509] = 10'd6;
  assign mem[2510] = 10'd6;
  assign mem[2511] = 10'd5;
  assign mem[2512] = 10'd4;
  assign mem[2513] = 10'd3;
  assign mem[2514] = 10'd2;
  assign mem[2515] = 10'd1;
  assign mem[2516] = 10'd2;
  assign mem[2517] = 10'd3;
  assign mem[2518] = 10'd4;
  assign mem[2519] = 10'd5;
  assign mem[2520] = 10'd5;
  assign mem[2521] = 10'd4;
  assign mem[2522] = 10'd3;
  assign mem[2523] = 10'd2;
  assign mem[2524] = 10'd1;
  assign mem[2525] = 10'd0;
  assign mem[2526] = 10'd1;
  assign mem[2527] = 10'd2;
  assign mem[2528] = 10'd3;
  assign mem[2529] = 10'd4;
  assign mem[2530] = 10'd6;
  assign mem[2531] = 10'd5;
  assign mem[2532] = 10'd4;
  assign mem[2533] = 10'd3;
  assign mem[2534] = 10'd2;
  assign mem[2535] = 10'd1;
  assign mem[2536] = 10'd2;
  assign mem[2537] = 10'd3;
  assign mem[2538] = 10'd4;
  assign mem[2539] = 10'd5;
  assign mem[2540] = 10'd7;
  assign mem[2541] = 10'd6;
  assign mem[2542] = 10'd5;
  assign mem[2543] = 10'd4;
  assign mem[2544] = 10'd3;
  assign mem[2545] = 10'd2;
  assign mem[2546] = 10'd3;
  assign mem[2547] = 10'd4;
  assign mem[2548] = 10'd5;
  assign mem[2549] = 10'd6;
  assign mem[2550] = 10'd8;
  assign mem[2551] = 10'd7;
  assign mem[2552] = 10'd6;
  assign mem[2553] = 10'd5;
  assign mem[2554] = 10'd4;
  assign mem[2555] = 10'd3;
  assign mem[2556] = 10'd4;
  assign mem[2557] = 10'd5;
  assign mem[2558] = 10'd6;
  assign mem[2559] = 10'd7;
  assign mem[2560] = 10'd9;
  assign mem[2561] = 10'd8;
  assign mem[2562] = 10'd7;
  assign mem[2563] = 10'd6;
  assign mem[2564] = 10'd5;
  assign mem[2565] = 10'd4;
  assign mem[2566] = 10'd5;
  assign mem[2567] = 10'd6;
  assign mem[2568] = 10'd7;
  assign mem[2569] = 10'd8;
  assign mem[2570] = 10'd10;
  assign mem[2571] = 10'd9;
  assign mem[2572] = 10'd8;
  assign mem[2573] = 10'd7;
  assign mem[2574] = 10'd6;
  assign mem[2575] = 10'd5;
  assign mem[2576] = 10'd6;
  assign mem[2577] = 10'd7;
  assign mem[2578] = 10'd8;
  assign mem[2579] = 10'd9;
  assign mem[2580] = 10'd11;
  assign mem[2581] = 10'd10;
  assign mem[2582] = 10'd9;
  assign mem[2583] = 10'd8;
  assign mem[2584] = 10'd7;
  assign mem[2585] = 10'd6;
  assign mem[2586] = 10'd7;
  assign mem[2587] = 10'd8;
  assign mem[2588] = 10'd9;
  assign mem[2589] = 10'd10;
  assign mem[2590] = 10'd12;
  assign mem[2591] = 10'd11;
  assign mem[2592] = 10'd10;
  assign mem[2593] = 10'd9;
  assign mem[2594] = 10'd8;
  assign mem[2595] = 10'd7;
  assign mem[2596] = 10'd8;
  assign mem[2597] = 10'd9;
  assign mem[2598] = 10'd10;
  assign mem[2599] = 10'd11;
  assign mem[2600] = 10'd8;
  assign mem[2601] = 10'd7;
  assign mem[2602] = 10'd6;
  assign mem[2603] = 10'd5;
  assign mem[2604] = 10'd4;
  assign mem[2605] = 10'd3;
  assign mem[2606] = 10'd2;
  assign mem[2607] = 10'd3;
  assign mem[2608] = 10'd4;
  assign mem[2609] = 10'd5;
  assign mem[2610] = 10'd7;
  assign mem[2611] = 10'd6;
  assign mem[2612] = 10'd5;
  assign mem[2613] = 10'd4;
  assign mem[2614] = 10'd3;
  assign mem[2615] = 10'd2;
  assign mem[2616] = 10'd1;
  assign mem[2617] = 10'd2;
  assign mem[2618] = 10'd3;
  assign mem[2619] = 10'd4;
  assign mem[2620] = 10'd6;
  assign mem[2621] = 10'd5;
  assign mem[2622] = 10'd4;
  assign mem[2623] = 10'd3;
  assign mem[2624] = 10'd2;
  assign mem[2625] = 10'd1;
  assign mem[2626] = 10'd0;
  assign mem[2627] = 10'd1;
  assign mem[2628] = 10'd2;
  assign mem[2629] = 10'd3;
  assign mem[2630] = 10'd7;
  assign mem[2631] = 10'd6;
  assign mem[2632] = 10'd5;
  assign mem[2633] = 10'd4;
  assign mem[2634] = 10'd3;
  assign mem[2635] = 10'd2;
  assign mem[2636] = 10'd1;
  assign mem[2637] = 10'd2;
  assign mem[2638] = 10'd3;
  assign mem[2639] = 10'd4;
  assign mem[2640] = 10'd8;
  assign mem[2641] = 10'd7;
  assign mem[2642] = 10'd6;
  assign mem[2643] = 10'd5;
  assign mem[2644] = 10'd4;
  assign mem[2645] = 10'd3;
  assign mem[2646] = 10'd2;
  assign mem[2647] = 10'd3;
  assign mem[2648] = 10'd4;
  assign mem[2649] = 10'd5;
  assign mem[2650] = 10'd9;
  assign mem[2651] = 10'd8;
  assign mem[2652] = 10'd7;
  assign mem[2653] = 10'd6;
  assign mem[2654] = 10'd5;
  assign mem[2655] = 10'd4;
  assign mem[2656] = 10'd3;
  assign mem[2657] = 10'd4;
  assign mem[2658] = 10'd5;
  assign mem[2659] = 10'd6;
  assign mem[2660] = 10'd10;
  assign mem[2661] = 10'd9;
  assign mem[2662] = 10'd8;
  assign mem[2663] = 10'd7;
  assign mem[2664] = 10'd6;
  assign mem[2665] = 10'd5;
  assign mem[2666] = 10'd4;
  assign mem[2667] = 10'd5;
  assign mem[2668] = 10'd6;
  assign mem[2669] = 10'd7;
  assign mem[2670] = 10'd11;
  assign mem[2671] = 10'd10;
  assign mem[2672] = 10'd9;
  assign mem[2673] = 10'd8;
  assign mem[2674] = 10'd7;
  assign mem[2675] = 10'd6;
  assign mem[2676] = 10'd5;
  assign mem[2677] = 10'd6;
  assign mem[2678] = 10'd7;
  assign mem[2679] = 10'd8;
  assign mem[2680] = 10'd12;
  assign mem[2681] = 10'd11;
  assign mem[2682] = 10'd10;
  assign mem[2683] = 10'd9;
  assign mem[2684] = 10'd8;
  assign mem[2685] = 10'd7;
  assign mem[2686] = 10'd6;
  assign mem[2687] = 10'd7;
  assign mem[2688] = 10'd8;
  assign mem[2689] = 10'd9;
  assign mem[2690] = 10'd13;
  assign mem[2691] = 10'd12;
  assign mem[2692] = 10'd11;
  assign mem[2693] = 10'd10;
  assign mem[2694] = 10'd9;
  assign mem[2695] = 10'd8;
  assign mem[2696] = 10'd7;
  assign mem[2697] = 10'd8;
  assign mem[2698] = 10'd9;
  assign mem[2699] = 10'd10;
  assign mem[2700] = 10'd9;
  assign mem[2701] = 10'd8;
  assign mem[2702] = 10'd7;
  assign mem[2703] = 10'd6;
  assign mem[2704] = 10'd5;
  assign mem[2705] = 10'd4;
  assign mem[2706] = 10'd3;
  assign mem[2707] = 10'd2;
  assign mem[2708] = 10'd3;
  assign mem[2709] = 10'd4;
  assign mem[2710] = 10'd8;
  assign mem[2711] = 10'd7;
  assign mem[2712] = 10'd6;
  assign mem[2713] = 10'd5;
  assign mem[2714] = 10'd4;
  assign mem[2715] = 10'd3;
  assign mem[2716] = 10'd2;
  assign mem[2717] = 10'd1;
  assign mem[2718] = 10'd2;
  assign mem[2719] = 10'd3;
  assign mem[2720] = 10'd7;
  assign mem[2721] = 10'd6;
  assign mem[2722] = 10'd5;
  assign mem[2723] = 10'd4;
  assign mem[2724] = 10'd3;
  assign mem[2725] = 10'd2;
  assign mem[2726] = 10'd1;
  assign mem[2727] = 10'd0;
  assign mem[2728] = 10'd1;
  assign mem[2729] = 10'd2;
  assign mem[2730] = 10'd8;
  assign mem[2731] = 10'd7;
  assign mem[2732] = 10'd6;
  assign mem[2733] = 10'd5;
  assign mem[2734] = 10'd4;
  assign mem[2735] = 10'd3;
  assign mem[2736] = 10'd2;
  assign mem[2737] = 10'd1;
  assign mem[2738] = 10'd2;
  assign mem[2739] = 10'd3;
  assign mem[2740] = 10'd9;
  assign mem[2741] = 10'd8;
  assign mem[2742] = 10'd7;
  assign mem[2743] = 10'd6;
  assign mem[2744] = 10'd5;
  assign mem[2745] = 10'd4;
  assign mem[2746] = 10'd3;
  assign mem[2747] = 10'd2;
  assign mem[2748] = 10'd3;
  assign mem[2749] = 10'd4;
  assign mem[2750] = 10'd10;
  assign mem[2751] = 10'd9;
  assign mem[2752] = 10'd8;
  assign mem[2753] = 10'd7;
  assign mem[2754] = 10'd6;
  assign mem[2755] = 10'd5;
  assign mem[2756] = 10'd4;
  assign mem[2757] = 10'd3;
  assign mem[2758] = 10'd4;
  assign mem[2759] = 10'd5;
  assign mem[2760] = 10'd11;
  assign mem[2761] = 10'd10;
  assign mem[2762] = 10'd9;
  assign mem[2763] = 10'd8;
  assign mem[2764] = 10'd7;
  assign mem[2765] = 10'd6;
  assign mem[2766] = 10'd5;
  assign mem[2767] = 10'd4;
  assign mem[2768] = 10'd5;
  assign mem[2769] = 10'd6;
  assign mem[2770] = 10'd12;
  assign mem[2771] = 10'd11;
  assign mem[2772] = 10'd10;
  assign mem[2773] = 10'd9;
  assign mem[2774] = 10'd8;
  assign mem[2775] = 10'd7;
  assign mem[2776] = 10'd6;
  assign mem[2777] = 10'd5;
  assign mem[2778] = 10'd6;
  assign mem[2779] = 10'd7;
  assign mem[2780] = 10'd13;
  assign mem[2781] = 10'd12;
  assign mem[2782] = 10'd11;
  assign mem[2783] = 10'd10;
  assign mem[2784] = 10'd9;
  assign mem[2785] = 10'd8;
  assign mem[2786] = 10'd7;
  assign mem[2787] = 10'd6;
  assign mem[2788] = 10'd7;
  assign mem[2789] = 10'd8;
  assign mem[2790] = 10'd14;
  assign mem[2791] = 10'd13;
  assign mem[2792] = 10'd12;
  assign mem[2793] = 10'd11;
  assign mem[2794] = 10'd10;
  assign mem[2795] = 10'd9;
  assign mem[2796] = 10'd8;
  assign mem[2797] = 10'd7;
  assign mem[2798] = 10'd8;
  assign mem[2799] = 10'd9;
  assign mem[2800] = 10'd10;
  assign mem[2801] = 10'd9;
  assign mem[2802] = 10'd8;
  assign mem[2803] = 10'd7;
  assign mem[2804] = 10'd6;
  assign mem[2805] = 10'd5;
  assign mem[2806] = 10'd4;
  assign mem[2807] = 10'd3;
  assign mem[2808] = 10'd2;
  assign mem[2809] = 10'd3;
  assign mem[2810] = 10'd9;
  assign mem[2811] = 10'd8;
  assign mem[2812] = 10'd7;
  assign mem[2813] = 10'd6;
  assign mem[2814] = 10'd5;
  assign mem[2815] = 10'd4;
  assign mem[2816] = 10'd3;
  assign mem[2817] = 10'd2;
  assign mem[2818] = 10'd1;
  assign mem[2819] = 10'd2;
  assign mem[2820] = 10'd8;
  assign mem[2821] = 10'd7;
  assign mem[2822] = 10'd6;
  assign mem[2823] = 10'd5;
  assign mem[2824] = 10'd4;
  assign mem[2825] = 10'd3;
  assign mem[2826] = 10'd2;
  assign mem[2827] = 10'd1;
  assign mem[2828] = 10'd0;
  assign mem[2829] = 10'd1;
  assign mem[2830] = 10'd9;
  assign mem[2831] = 10'd8;
  assign mem[2832] = 10'd7;
  assign mem[2833] = 10'd6;
  assign mem[2834] = 10'd5;
  assign mem[2835] = 10'd4;
  assign mem[2836] = 10'd3;
  assign mem[2837] = 10'd2;
  assign mem[2838] = 10'd1;
  assign mem[2839] = 10'd2;
  assign mem[2840] = 10'd10;
  assign mem[2841] = 10'd9;
  assign mem[2842] = 10'd8;
  assign mem[2843] = 10'd7;
  assign mem[2844] = 10'd6;
  assign mem[2845] = 10'd5;
  assign mem[2846] = 10'd4;
  assign mem[2847] = 10'd3;
  assign mem[2848] = 10'd2;
  assign mem[2849] = 10'd3;
  assign mem[2850] = 10'd11;
  assign mem[2851] = 10'd10;
  assign mem[2852] = 10'd9;
  assign mem[2853] = 10'd8;
  assign mem[2854] = 10'd7;
  assign mem[2855] = 10'd6;
  assign mem[2856] = 10'd5;
  assign mem[2857] = 10'd4;
  assign mem[2858] = 10'd3;
  assign mem[2859] = 10'd4;
  assign mem[2860] = 10'd12;
  assign mem[2861] = 10'd11;
  assign mem[2862] = 10'd10;
  assign mem[2863] = 10'd9;
  assign mem[2864] = 10'd8;
  assign mem[2865] = 10'd7;
  assign mem[2866] = 10'd6;
  assign mem[2867] = 10'd5;
  assign mem[2868] = 10'd4;
  assign mem[2869] = 10'd5;
  assign mem[2870] = 10'd13;
  assign mem[2871] = 10'd12;
  assign mem[2872] = 10'd11;
  assign mem[2873] = 10'd10;
  assign mem[2874] = 10'd9;
  assign mem[2875] = 10'd8;
  assign mem[2876] = 10'd7;
  assign mem[2877] = 10'd6;
  assign mem[2878] = 10'd5;
  assign mem[2879] = 10'd6;
  assign mem[2880] = 10'd14;
  assign mem[2881] = 10'd13;
  assign mem[2882] = 10'd12;
  assign mem[2883] = 10'd11;
  assign mem[2884] = 10'd10;
  assign mem[2885] = 10'd9;
  assign mem[2886] = 10'd8;
  assign mem[2887] = 10'd7;
  assign mem[2888] = 10'd6;
  assign mem[2889] = 10'd7;
  assign mem[2890] = 10'd15;
  assign mem[2891] = 10'd14;
  assign mem[2892] = 10'd13;
  assign mem[2893] = 10'd12;
  assign mem[2894] = 10'd11;
  assign mem[2895] = 10'd10;
  assign mem[2896] = 10'd9;
  assign mem[2897] = 10'd8;
  assign mem[2898] = 10'd7;
  assign mem[2899] = 10'd8;
  assign mem[2900] = 10'd11;
  assign mem[2901] = 10'd10;
  assign mem[2902] = 10'd9;
  assign mem[2903] = 10'd8;
  assign mem[2904] = 10'd7;
  assign mem[2905] = 10'd6;
  assign mem[2906] = 10'd5;
  assign mem[2907] = 10'd4;
  assign mem[2908] = 10'd3;
  assign mem[2909] = 10'd2;
  assign mem[2910] = 10'd10;
  assign mem[2911] = 10'd9;
  assign mem[2912] = 10'd8;
  assign mem[2913] = 10'd7;
  assign mem[2914] = 10'd6;
  assign mem[2915] = 10'd5;
  assign mem[2916] = 10'd4;
  assign mem[2917] = 10'd3;
  assign mem[2918] = 10'd2;
  assign mem[2919] = 10'd1;
  assign mem[2920] = 10'd9;
  assign mem[2921] = 10'd8;
  assign mem[2922] = 10'd7;
  assign mem[2923] = 10'd6;
  assign mem[2924] = 10'd5;
  assign mem[2925] = 10'd4;
  assign mem[2926] = 10'd3;
  assign mem[2927] = 10'd2;
  assign mem[2928] = 10'd1;
  assign mem[2929] = 10'd0;
  assign mem[2930] = 10'd10;
  assign mem[2931] = 10'd9;
  assign mem[2932] = 10'd8;
  assign mem[2933] = 10'd7;
  assign mem[2934] = 10'd6;
  assign mem[2935] = 10'd5;
  assign mem[2936] = 10'd4;
  assign mem[2937] = 10'd3;
  assign mem[2938] = 10'd2;
  assign mem[2939] = 10'd1;
  assign mem[2940] = 10'd11;
  assign mem[2941] = 10'd10;
  assign mem[2942] = 10'd9;
  assign mem[2943] = 10'd8;
  assign mem[2944] = 10'd7;
  assign mem[2945] = 10'd6;
  assign mem[2946] = 10'd5;
  assign mem[2947] = 10'd4;
  assign mem[2948] = 10'd3;
  assign mem[2949] = 10'd2;
  assign mem[2950] = 10'd12;
  assign mem[2951] = 10'd11;
  assign mem[2952] = 10'd10;
  assign mem[2953] = 10'd9;
  assign mem[2954] = 10'd8;
  assign mem[2955] = 10'd7;
  assign mem[2956] = 10'd6;
  assign mem[2957] = 10'd5;
  assign mem[2958] = 10'd4;
  assign mem[2959] = 10'd3;
  assign mem[2960] = 10'd13;
  assign mem[2961] = 10'd12;
  assign mem[2962] = 10'd11;
  assign mem[2963] = 10'd10;
  assign mem[2964] = 10'd9;
  assign mem[2965] = 10'd8;
  assign mem[2966] = 10'd7;
  assign mem[2967] = 10'd6;
  assign mem[2968] = 10'd5;
  assign mem[2969] = 10'd4;
  assign mem[2970] = 10'd14;
  assign mem[2971] = 10'd13;
  assign mem[2972] = 10'd12;
  assign mem[2973] = 10'd11;
  assign mem[2974] = 10'd10;
  assign mem[2975] = 10'd9;
  assign mem[2976] = 10'd8;
  assign mem[2977] = 10'd7;
  assign mem[2978] = 10'd6;
  assign mem[2979] = 10'd5;
  assign mem[2980] = 10'd15;
  assign mem[2981] = 10'd14;
  assign mem[2982] = 10'd13;
  assign mem[2983] = 10'd12;
  assign mem[2984] = 10'd11;
  assign mem[2985] = 10'd10;
  assign mem[2986] = 10'd9;
  assign mem[2987] = 10'd8;
  assign mem[2988] = 10'd7;
  assign mem[2989] = 10'd6;
  assign mem[2990] = 10'd16;
  assign mem[2991] = 10'd15;
  assign mem[2992] = 10'd14;
  assign mem[2993] = 10'd13;
  assign mem[2994] = 10'd12;
  assign mem[2995] = 10'd11;
  assign mem[2996] = 10'd10;
  assign mem[2997] = 10'd9;
  assign mem[2998] = 10'd8;
  assign mem[2999] = 10'd7;
  assign mem[3000] = 10'd3;
  assign mem[3001] = 10'd4;
  assign mem[3002] = 10'd5;
  assign mem[3003] = 10'd6;
  assign mem[3004] = 10'd7;
  assign mem[3005] = 10'd8;
  assign mem[3006] = 10'd9;
  assign mem[3007] = 10'd10;
  assign mem[3008] = 10'd11;
  assign mem[3009] = 10'd12;
  assign mem[3010] = 10'd2;
  assign mem[3011] = 10'd3;
  assign mem[3012] = 10'd4;
  assign mem[3013] = 10'd5;
  assign mem[3014] = 10'd6;
  assign mem[3015] = 10'd7;
  assign mem[3016] = 10'd8;
  assign mem[3017] = 10'd9;
  assign mem[3018] = 10'd10;
  assign mem[3019] = 10'd11;
  assign mem[3020] = 10'd1;
  assign mem[3021] = 10'd2;
  assign mem[3022] = 10'd3;
  assign mem[3023] = 10'd4;
  assign mem[3024] = 10'd5;
  assign mem[3025] = 10'd6;
  assign mem[3026] = 10'd7;
  assign mem[3027] = 10'd8;
  assign mem[3028] = 10'd9;
  assign mem[3029] = 10'd10;
  assign mem[3030] = 10'd0;
  assign mem[3031] = 10'd1;
  assign mem[3032] = 10'd2;
  assign mem[3033] = 10'd3;
  assign mem[3034] = 10'd4;
  assign mem[3035] = 10'd5;
  assign mem[3036] = 10'd6;
  assign mem[3037] = 10'd7;
  assign mem[3038] = 10'd8;
  assign mem[3039] = 10'd9;
  assign mem[3040] = 10'd1;
  assign mem[3041] = 10'd2;
  assign mem[3042] = 10'd3;
  assign mem[3043] = 10'd4;
  assign mem[3044] = 10'd5;
  assign mem[3045] = 10'd6;
  assign mem[3046] = 10'd7;
  assign mem[3047] = 10'd8;
  assign mem[3048] = 10'd9;
  assign mem[3049] = 10'd10;
  assign mem[3050] = 10'd2;
  assign mem[3051] = 10'd3;
  assign mem[3052] = 10'd4;
  assign mem[3053] = 10'd5;
  assign mem[3054] = 10'd6;
  assign mem[3055] = 10'd7;
  assign mem[3056] = 10'd8;
  assign mem[3057] = 10'd9;
  assign mem[3058] = 10'd10;
  assign mem[3059] = 10'd11;
  assign mem[3060] = 10'd3;
  assign mem[3061] = 10'd4;
  assign mem[3062] = 10'd5;
  assign mem[3063] = 10'd6;
  assign mem[3064] = 10'd7;
  assign mem[3065] = 10'd8;
  assign mem[3066] = 10'd9;
  assign mem[3067] = 10'd10;
  assign mem[3068] = 10'd11;
  assign mem[3069] = 10'd12;
  assign mem[3070] = 10'd4;
  assign mem[3071] = 10'd5;
  assign mem[3072] = 10'd6;
  assign mem[3073] = 10'd7;
  assign mem[3074] = 10'd8;
  assign mem[3075] = 10'd9;
  assign mem[3076] = 10'd10;
  assign mem[3077] = 10'd11;
  assign mem[3078] = 10'd12;
  assign mem[3079] = 10'd13;
  assign mem[3080] = 10'd5;
  assign mem[3081] = 10'd6;
  assign mem[3082] = 10'd7;
  assign mem[3083] = 10'd8;
  assign mem[3084] = 10'd9;
  assign mem[3085] = 10'd10;
  assign mem[3086] = 10'd11;
  assign mem[3087] = 10'd12;
  assign mem[3088] = 10'd13;
  assign mem[3089] = 10'd14;
  assign mem[3090] = 10'd6;
  assign mem[3091] = 10'd7;
  assign mem[3092] = 10'd8;
  assign mem[3093] = 10'd9;
  assign mem[3094] = 10'd10;
  assign mem[3095] = 10'd11;
  assign mem[3096] = 10'd12;
  assign mem[3097] = 10'd13;
  assign mem[3098] = 10'd14;
  assign mem[3099] = 10'd15;
  assign mem[3100] = 10'd4;
  assign mem[3101] = 10'd3;
  assign mem[3102] = 10'd4;
  assign mem[3103] = 10'd5;
  assign mem[3104] = 10'd6;
  assign mem[3105] = 10'd7;
  assign mem[3106] = 10'd8;
  assign mem[3107] = 10'd9;
  assign mem[3108] = 10'd10;
  assign mem[3109] = 10'd11;
  assign mem[3110] = 10'd3;
  assign mem[3111] = 10'd2;
  assign mem[3112] = 10'd3;
  assign mem[3113] = 10'd4;
  assign mem[3114] = 10'd5;
  assign mem[3115] = 10'd6;
  assign mem[3116] = 10'd7;
  assign mem[3117] = 10'd8;
  assign mem[3118] = 10'd9;
  assign mem[3119] = 10'd10;
  assign mem[3120] = 10'd2;
  assign mem[3121] = 10'd1;
  assign mem[3122] = 10'd2;
  assign mem[3123] = 10'd3;
  assign mem[3124] = 10'd4;
  assign mem[3125] = 10'd5;
  assign mem[3126] = 10'd6;
  assign mem[3127] = 10'd7;
  assign mem[3128] = 10'd8;
  assign mem[3129] = 10'd9;
  assign mem[3130] = 10'd1;
  assign mem[3131] = 10'd0;
  assign mem[3132] = 10'd1;
  assign mem[3133] = 10'd2;
  assign mem[3134] = 10'd3;
  assign mem[3135] = 10'd4;
  assign mem[3136] = 10'd5;
  assign mem[3137] = 10'd6;
  assign mem[3138] = 10'd7;
  assign mem[3139] = 10'd8;
  assign mem[3140] = 10'd2;
  assign mem[3141] = 10'd1;
  assign mem[3142] = 10'd2;
  assign mem[3143] = 10'd3;
  assign mem[3144] = 10'd4;
  assign mem[3145] = 10'd5;
  assign mem[3146] = 10'd6;
  assign mem[3147] = 10'd7;
  assign mem[3148] = 10'd8;
  assign mem[3149] = 10'd9;
  assign mem[3150] = 10'd3;
  assign mem[3151] = 10'd2;
  assign mem[3152] = 10'd3;
  assign mem[3153] = 10'd4;
  assign mem[3154] = 10'd5;
  assign mem[3155] = 10'd6;
  assign mem[3156] = 10'd7;
  assign mem[3157] = 10'd8;
  assign mem[3158] = 10'd9;
  assign mem[3159] = 10'd10;
  assign mem[3160] = 10'd4;
  assign mem[3161] = 10'd3;
  assign mem[3162] = 10'd4;
  assign mem[3163] = 10'd5;
  assign mem[3164] = 10'd6;
  assign mem[3165] = 10'd7;
  assign mem[3166] = 10'd8;
  assign mem[3167] = 10'd9;
  assign mem[3168] = 10'd10;
  assign mem[3169] = 10'd11;
  assign mem[3170] = 10'd5;
  assign mem[3171] = 10'd4;
  assign mem[3172] = 10'd5;
  assign mem[3173] = 10'd6;
  assign mem[3174] = 10'd7;
  assign mem[3175] = 10'd8;
  assign mem[3176] = 10'd9;
  assign mem[3177] = 10'd10;
  assign mem[3178] = 10'd11;
  assign mem[3179] = 10'd12;
  assign mem[3180] = 10'd6;
  assign mem[3181] = 10'd5;
  assign mem[3182] = 10'd6;
  assign mem[3183] = 10'd7;
  assign mem[3184] = 10'd8;
  assign mem[3185] = 10'd9;
  assign mem[3186] = 10'd10;
  assign mem[3187] = 10'd11;
  assign mem[3188] = 10'd12;
  assign mem[3189] = 10'd13;
  assign mem[3190] = 10'd7;
  assign mem[3191] = 10'd6;
  assign mem[3192] = 10'd7;
  assign mem[3193] = 10'd8;
  assign mem[3194] = 10'd9;
  assign mem[3195] = 10'd10;
  assign mem[3196] = 10'd11;
  assign mem[3197] = 10'd12;
  assign mem[3198] = 10'd13;
  assign mem[3199] = 10'd14;
  assign mem[3200] = 10'd5;
  assign mem[3201] = 10'd4;
  assign mem[3202] = 10'd3;
  assign mem[3203] = 10'd4;
  assign mem[3204] = 10'd5;
  assign mem[3205] = 10'd6;
  assign mem[3206] = 10'd7;
  assign mem[3207] = 10'd8;
  assign mem[3208] = 10'd9;
  assign mem[3209] = 10'd10;
  assign mem[3210] = 10'd4;
  assign mem[3211] = 10'd3;
  assign mem[3212] = 10'd2;
  assign mem[3213] = 10'd3;
  assign mem[3214] = 10'd4;
  assign mem[3215] = 10'd5;
  assign mem[3216] = 10'd6;
  assign mem[3217] = 10'd7;
  assign mem[3218] = 10'd8;
  assign mem[3219] = 10'd9;
  assign mem[3220] = 10'd3;
  assign mem[3221] = 10'd2;
  assign mem[3222] = 10'd1;
  assign mem[3223] = 10'd2;
  assign mem[3224] = 10'd3;
  assign mem[3225] = 10'd4;
  assign mem[3226] = 10'd5;
  assign mem[3227] = 10'd6;
  assign mem[3228] = 10'd7;
  assign mem[3229] = 10'd8;
  assign mem[3230] = 10'd2;
  assign mem[3231] = 10'd1;
  assign mem[3232] = 10'd0;
  assign mem[3233] = 10'd1;
  assign mem[3234] = 10'd2;
  assign mem[3235] = 10'd3;
  assign mem[3236] = 10'd4;
  assign mem[3237] = 10'd5;
  assign mem[3238] = 10'd6;
  assign mem[3239] = 10'd7;
  assign mem[3240] = 10'd3;
  assign mem[3241] = 10'd2;
  assign mem[3242] = 10'd1;
  assign mem[3243] = 10'd2;
  assign mem[3244] = 10'd3;
  assign mem[3245] = 10'd4;
  assign mem[3246] = 10'd5;
  assign mem[3247] = 10'd6;
  assign mem[3248] = 10'd7;
  assign mem[3249] = 10'd8;
  assign mem[3250] = 10'd4;
  assign mem[3251] = 10'd3;
  assign mem[3252] = 10'd2;
  assign mem[3253] = 10'd3;
  assign mem[3254] = 10'd4;
  assign mem[3255] = 10'd5;
  assign mem[3256] = 10'd6;
  assign mem[3257] = 10'd7;
  assign mem[3258] = 10'd8;
  assign mem[3259] = 10'd9;
  assign mem[3260] = 10'd5;
  assign mem[3261] = 10'd4;
  assign mem[3262] = 10'd3;
  assign mem[3263] = 10'd4;
  assign mem[3264] = 10'd5;
  assign mem[3265] = 10'd6;
  assign mem[3266] = 10'd7;
  assign mem[3267] = 10'd8;
  assign mem[3268] = 10'd9;
  assign mem[3269] = 10'd10;
  assign mem[3270] = 10'd6;
  assign mem[3271] = 10'd5;
  assign mem[3272] = 10'd4;
  assign mem[3273] = 10'd5;
  assign mem[3274] = 10'd6;
  assign mem[3275] = 10'd7;
  assign mem[3276] = 10'd8;
  assign mem[3277] = 10'd9;
  assign mem[3278] = 10'd10;
  assign mem[3279] = 10'd11;
  assign mem[3280] = 10'd7;
  assign mem[3281] = 10'd6;
  assign mem[3282] = 10'd5;
  assign mem[3283] = 10'd6;
  assign mem[3284] = 10'd7;
  assign mem[3285] = 10'd8;
  assign mem[3286] = 10'd9;
  assign mem[3287] = 10'd10;
  assign mem[3288] = 10'd11;
  assign mem[3289] = 10'd12;
  assign mem[3290] = 10'd8;
  assign mem[3291] = 10'd7;
  assign mem[3292] = 10'd6;
  assign mem[3293] = 10'd7;
  assign mem[3294] = 10'd8;
  assign mem[3295] = 10'd9;
  assign mem[3296] = 10'd10;
  assign mem[3297] = 10'd11;
  assign mem[3298] = 10'd12;
  assign mem[3299] = 10'd13;
  assign mem[3300] = 10'd6;
  assign mem[3301] = 10'd5;
  assign mem[3302] = 10'd4;
  assign mem[3303] = 10'd3;
  assign mem[3304] = 10'd4;
  assign mem[3305] = 10'd5;
  assign mem[3306] = 10'd6;
  assign mem[3307] = 10'd7;
  assign mem[3308] = 10'd8;
  assign mem[3309] = 10'd9;
  assign mem[3310] = 10'd5;
  assign mem[3311] = 10'd4;
  assign mem[3312] = 10'd3;
  assign mem[3313] = 10'd2;
  assign mem[3314] = 10'd3;
  assign mem[3315] = 10'd4;
  assign mem[3316] = 10'd5;
  assign mem[3317] = 10'd6;
  assign mem[3318] = 10'd7;
  assign mem[3319] = 10'd8;
  assign mem[3320] = 10'd4;
  assign mem[3321] = 10'd3;
  assign mem[3322] = 10'd2;
  assign mem[3323] = 10'd1;
  assign mem[3324] = 10'd2;
  assign mem[3325] = 10'd3;
  assign mem[3326] = 10'd4;
  assign mem[3327] = 10'd5;
  assign mem[3328] = 10'd6;
  assign mem[3329] = 10'd7;
  assign mem[3330] = 10'd3;
  assign mem[3331] = 10'd2;
  assign mem[3332] = 10'd1;
  assign mem[3333] = 10'd0;
  assign mem[3334] = 10'd1;
  assign mem[3335] = 10'd2;
  assign mem[3336] = 10'd3;
  assign mem[3337] = 10'd4;
  assign mem[3338] = 10'd5;
  assign mem[3339] = 10'd6;
  assign mem[3340] = 10'd4;
  assign mem[3341] = 10'd3;
  assign mem[3342] = 10'd2;
  assign mem[3343] = 10'd1;
  assign mem[3344] = 10'd2;
  assign mem[3345] = 10'd3;
  assign mem[3346] = 10'd4;
  assign mem[3347] = 10'd5;
  assign mem[3348] = 10'd6;
  assign mem[3349] = 10'd7;
  assign mem[3350] = 10'd5;
  assign mem[3351] = 10'd4;
  assign mem[3352] = 10'd3;
  assign mem[3353] = 10'd2;
  assign mem[3354] = 10'd3;
  assign mem[3355] = 10'd4;
  assign mem[3356] = 10'd5;
  assign mem[3357] = 10'd6;
  assign mem[3358] = 10'd7;
  assign mem[3359] = 10'd8;
  assign mem[3360] = 10'd6;
  assign mem[3361] = 10'd5;
  assign mem[3362] = 10'd4;
  assign mem[3363] = 10'd3;
  assign mem[3364] = 10'd4;
  assign mem[3365] = 10'd5;
  assign mem[3366] = 10'd6;
  assign mem[3367] = 10'd7;
  assign mem[3368] = 10'd8;
  assign mem[3369] = 10'd9;
  assign mem[3370] = 10'd7;
  assign mem[3371] = 10'd6;
  assign mem[3372] = 10'd5;
  assign mem[3373] = 10'd4;
  assign mem[3374] = 10'd5;
  assign mem[3375] = 10'd6;
  assign mem[3376] = 10'd7;
  assign mem[3377] = 10'd8;
  assign mem[3378] = 10'd9;
  assign mem[3379] = 10'd10;
  assign mem[3380] = 10'd8;
  assign mem[3381] = 10'd7;
  assign mem[3382] = 10'd6;
  assign mem[3383] = 10'd5;
  assign mem[3384] = 10'd6;
  assign mem[3385] = 10'd7;
  assign mem[3386] = 10'd8;
  assign mem[3387] = 10'd9;
  assign mem[3388] = 10'd10;
  assign mem[3389] = 10'd11;
  assign mem[3390] = 10'd9;
  assign mem[3391] = 10'd8;
  assign mem[3392] = 10'd7;
  assign mem[3393] = 10'd6;
  assign mem[3394] = 10'd7;
  assign mem[3395] = 10'd8;
  assign mem[3396] = 10'd9;
  assign mem[3397] = 10'd10;
  assign mem[3398] = 10'd11;
  assign mem[3399] = 10'd12;
  assign mem[3400] = 10'd7;
  assign mem[3401] = 10'd6;
  assign mem[3402] = 10'd5;
  assign mem[3403] = 10'd4;
  assign mem[3404] = 10'd3;
  assign mem[3405] = 10'd4;
  assign mem[3406] = 10'd5;
  assign mem[3407] = 10'd6;
  assign mem[3408] = 10'd7;
  assign mem[3409] = 10'd8;
  assign mem[3410] = 10'd6;
  assign mem[3411] = 10'd5;
  assign mem[3412] = 10'd4;
  assign mem[3413] = 10'd3;
  assign mem[3414] = 10'd2;
  assign mem[3415] = 10'd3;
  assign mem[3416] = 10'd4;
  assign mem[3417] = 10'd5;
  assign mem[3418] = 10'd6;
  assign mem[3419] = 10'd7;
  assign mem[3420] = 10'd5;
  assign mem[3421] = 10'd4;
  assign mem[3422] = 10'd3;
  assign mem[3423] = 10'd2;
  assign mem[3424] = 10'd1;
  assign mem[3425] = 10'd2;
  assign mem[3426] = 10'd3;
  assign mem[3427] = 10'd4;
  assign mem[3428] = 10'd5;
  assign mem[3429] = 10'd6;
  assign mem[3430] = 10'd4;
  assign mem[3431] = 10'd3;
  assign mem[3432] = 10'd2;
  assign mem[3433] = 10'd1;
  assign mem[3434] = 10'd0;
  assign mem[3435] = 10'd1;
  assign mem[3436] = 10'd2;
  assign mem[3437] = 10'd3;
  assign mem[3438] = 10'd4;
  assign mem[3439] = 10'd5;
  assign mem[3440] = 10'd5;
  assign mem[3441] = 10'd4;
  assign mem[3442] = 10'd3;
  assign mem[3443] = 10'd2;
  assign mem[3444] = 10'd1;
  assign mem[3445] = 10'd2;
  assign mem[3446] = 10'd3;
  assign mem[3447] = 10'd4;
  assign mem[3448] = 10'd5;
  assign mem[3449] = 10'd6;
  assign mem[3450] = 10'd6;
  assign mem[3451] = 10'd5;
  assign mem[3452] = 10'd4;
  assign mem[3453] = 10'd3;
  assign mem[3454] = 10'd2;
  assign mem[3455] = 10'd3;
  assign mem[3456] = 10'd4;
  assign mem[3457] = 10'd5;
  assign mem[3458] = 10'd6;
  assign mem[3459] = 10'd7;
  assign mem[3460] = 10'd7;
  assign mem[3461] = 10'd6;
  assign mem[3462] = 10'd5;
  assign mem[3463] = 10'd4;
  assign mem[3464] = 10'd3;
  assign mem[3465] = 10'd4;
  assign mem[3466] = 10'd5;
  assign mem[3467] = 10'd6;
  assign mem[3468] = 10'd7;
  assign mem[3469] = 10'd8;
  assign mem[3470] = 10'd8;
  assign mem[3471] = 10'd7;
  assign mem[3472] = 10'd6;
  assign mem[3473] = 10'd5;
  assign mem[3474] = 10'd4;
  assign mem[3475] = 10'd5;
  assign mem[3476] = 10'd6;
  assign mem[3477] = 10'd7;
  assign mem[3478] = 10'd8;
  assign mem[3479] = 10'd9;
  assign mem[3480] = 10'd9;
  assign mem[3481] = 10'd8;
  assign mem[3482] = 10'd7;
  assign mem[3483] = 10'd6;
  assign mem[3484] = 10'd5;
  assign mem[3485] = 10'd6;
  assign mem[3486] = 10'd7;
  assign mem[3487] = 10'd8;
  assign mem[3488] = 10'd9;
  assign mem[3489] = 10'd10;
  assign mem[3490] = 10'd10;
  assign mem[3491] = 10'd9;
  assign mem[3492] = 10'd8;
  assign mem[3493] = 10'd7;
  assign mem[3494] = 10'd6;
  assign mem[3495] = 10'd7;
  assign mem[3496] = 10'd8;
  assign mem[3497] = 10'd9;
  assign mem[3498] = 10'd10;
  assign mem[3499] = 10'd11;
  assign mem[3500] = 10'd8;
  assign mem[3501] = 10'd7;
  assign mem[3502] = 10'd6;
  assign mem[3503] = 10'd5;
  assign mem[3504] = 10'd4;
  assign mem[3505] = 10'd3;
  assign mem[3506] = 10'd4;
  assign mem[3507] = 10'd5;
  assign mem[3508] = 10'd6;
  assign mem[3509] = 10'd7;
  assign mem[3510] = 10'd7;
  assign mem[3511] = 10'd6;
  assign mem[3512] = 10'd5;
  assign mem[3513] = 10'd4;
  assign mem[3514] = 10'd3;
  assign mem[3515] = 10'd2;
  assign mem[3516] = 10'd3;
  assign mem[3517] = 10'd4;
  assign mem[3518] = 10'd5;
  assign mem[3519] = 10'd6;
  assign mem[3520] = 10'd6;
  assign mem[3521] = 10'd5;
  assign mem[3522] = 10'd4;
  assign mem[3523] = 10'd3;
  assign mem[3524] = 10'd2;
  assign mem[3525] = 10'd1;
  assign mem[3526] = 10'd2;
  assign mem[3527] = 10'd3;
  assign mem[3528] = 10'd4;
  assign mem[3529] = 10'd5;
  assign mem[3530] = 10'd5;
  assign mem[3531] = 10'd4;
  assign mem[3532] = 10'd3;
  assign mem[3533] = 10'd2;
  assign mem[3534] = 10'd1;
  assign mem[3535] = 10'd0;
  assign mem[3536] = 10'd1;
  assign mem[3537] = 10'd2;
  assign mem[3538] = 10'd3;
  assign mem[3539] = 10'd4;
  assign mem[3540] = 10'd6;
  assign mem[3541] = 10'd5;
  assign mem[3542] = 10'd4;
  assign mem[3543] = 10'd3;
  assign mem[3544] = 10'd2;
  assign mem[3545] = 10'd1;
  assign mem[3546] = 10'd2;
  assign mem[3547] = 10'd3;
  assign mem[3548] = 10'd4;
  assign mem[3549] = 10'd5;
  assign mem[3550] = 10'd7;
  assign mem[3551] = 10'd6;
  assign mem[3552] = 10'd5;
  assign mem[3553] = 10'd4;
  assign mem[3554] = 10'd3;
  assign mem[3555] = 10'd2;
  assign mem[3556] = 10'd3;
  assign mem[3557] = 10'd4;
  assign mem[3558] = 10'd5;
  assign mem[3559] = 10'd6;
  assign mem[3560] = 10'd8;
  assign mem[3561] = 10'd7;
  assign mem[3562] = 10'd6;
  assign mem[3563] = 10'd5;
  assign mem[3564] = 10'd4;
  assign mem[3565] = 10'd3;
  assign mem[3566] = 10'd4;
  assign mem[3567] = 10'd5;
  assign mem[3568] = 10'd6;
  assign mem[3569] = 10'd7;
  assign mem[3570] = 10'd9;
  assign mem[3571] = 10'd8;
  assign mem[3572] = 10'd7;
  assign mem[3573] = 10'd6;
  assign mem[3574] = 10'd5;
  assign mem[3575] = 10'd4;
  assign mem[3576] = 10'd5;
  assign mem[3577] = 10'd6;
  assign mem[3578] = 10'd7;
  assign mem[3579] = 10'd8;
  assign mem[3580] = 10'd10;
  assign mem[3581] = 10'd9;
  assign mem[3582] = 10'd8;
  assign mem[3583] = 10'd7;
  assign mem[3584] = 10'd6;
  assign mem[3585] = 10'd5;
  assign mem[3586] = 10'd6;
  assign mem[3587] = 10'd7;
  assign mem[3588] = 10'd8;
  assign mem[3589] = 10'd9;
  assign mem[3590] = 10'd11;
  assign mem[3591] = 10'd10;
  assign mem[3592] = 10'd9;
  assign mem[3593] = 10'd8;
  assign mem[3594] = 10'd7;
  assign mem[3595] = 10'd6;
  assign mem[3596] = 10'd7;
  assign mem[3597] = 10'd8;
  assign mem[3598] = 10'd9;
  assign mem[3599] = 10'd10;
  assign mem[3600] = 10'd9;
  assign mem[3601] = 10'd8;
  assign mem[3602] = 10'd7;
  assign mem[3603] = 10'd6;
  assign mem[3604] = 10'd5;
  assign mem[3605] = 10'd4;
  assign mem[3606] = 10'd3;
  assign mem[3607] = 10'd4;
  assign mem[3608] = 10'd5;
  assign mem[3609] = 10'd6;
  assign mem[3610] = 10'd8;
  assign mem[3611] = 10'd7;
  assign mem[3612] = 10'd6;
  assign mem[3613] = 10'd5;
  assign mem[3614] = 10'd4;
  assign mem[3615] = 10'd3;
  assign mem[3616] = 10'd2;
  assign mem[3617] = 10'd3;
  assign mem[3618] = 10'd4;
  assign mem[3619] = 10'd5;
  assign mem[3620] = 10'd7;
  assign mem[3621] = 10'd6;
  assign mem[3622] = 10'd5;
  assign mem[3623] = 10'd4;
  assign mem[3624] = 10'd3;
  assign mem[3625] = 10'd2;
  assign mem[3626] = 10'd1;
  assign mem[3627] = 10'd2;
  assign mem[3628] = 10'd3;
  assign mem[3629] = 10'd4;
  assign mem[3630] = 10'd6;
  assign mem[3631] = 10'd5;
  assign mem[3632] = 10'd4;
  assign mem[3633] = 10'd3;
  assign mem[3634] = 10'd2;
  assign mem[3635] = 10'd1;
  assign mem[3636] = 10'd0;
  assign mem[3637] = 10'd1;
  assign mem[3638] = 10'd2;
  assign mem[3639] = 10'd3;
  assign mem[3640] = 10'd7;
  assign mem[3641] = 10'd6;
  assign mem[3642] = 10'd5;
  assign mem[3643] = 10'd4;
  assign mem[3644] = 10'd3;
  assign mem[3645] = 10'd2;
  assign mem[3646] = 10'd1;
  assign mem[3647] = 10'd2;
  assign mem[3648] = 10'd3;
  assign mem[3649] = 10'd4;
  assign mem[3650] = 10'd8;
  assign mem[3651] = 10'd7;
  assign mem[3652] = 10'd6;
  assign mem[3653] = 10'd5;
  assign mem[3654] = 10'd4;
  assign mem[3655] = 10'd3;
  assign mem[3656] = 10'd2;
  assign mem[3657] = 10'd3;
  assign mem[3658] = 10'd4;
  assign mem[3659] = 10'd5;
  assign mem[3660] = 10'd9;
  assign mem[3661] = 10'd8;
  assign mem[3662] = 10'd7;
  assign mem[3663] = 10'd6;
  assign mem[3664] = 10'd5;
  assign mem[3665] = 10'd4;
  assign mem[3666] = 10'd3;
  assign mem[3667] = 10'd4;
  assign mem[3668] = 10'd5;
  assign mem[3669] = 10'd6;
  assign mem[3670] = 10'd10;
  assign mem[3671] = 10'd9;
  assign mem[3672] = 10'd8;
  assign mem[3673] = 10'd7;
  assign mem[3674] = 10'd6;
  assign mem[3675] = 10'd5;
  assign mem[3676] = 10'd4;
  assign mem[3677] = 10'd5;
  assign mem[3678] = 10'd6;
  assign mem[3679] = 10'd7;
  assign mem[3680] = 10'd11;
  assign mem[3681] = 10'd10;
  assign mem[3682] = 10'd9;
  assign mem[3683] = 10'd8;
  assign mem[3684] = 10'd7;
  assign mem[3685] = 10'd6;
  assign mem[3686] = 10'd5;
  assign mem[3687] = 10'd6;
  assign mem[3688] = 10'd7;
  assign mem[3689] = 10'd8;
  assign mem[3690] = 10'd12;
  assign mem[3691] = 10'd11;
  assign mem[3692] = 10'd10;
  assign mem[3693] = 10'd9;
  assign mem[3694] = 10'd8;
  assign mem[3695] = 10'd7;
  assign mem[3696] = 10'd6;
  assign mem[3697] = 10'd7;
  assign mem[3698] = 10'd8;
  assign mem[3699] = 10'd9;
  assign mem[3700] = 10'd10;
  assign mem[3701] = 10'd9;
  assign mem[3702] = 10'd8;
  assign mem[3703] = 10'd7;
  assign mem[3704] = 10'd6;
  assign mem[3705] = 10'd5;
  assign mem[3706] = 10'd4;
  assign mem[3707] = 10'd3;
  assign mem[3708] = 10'd4;
  assign mem[3709] = 10'd5;
  assign mem[3710] = 10'd9;
  assign mem[3711] = 10'd8;
  assign mem[3712] = 10'd7;
  assign mem[3713] = 10'd6;
  assign mem[3714] = 10'd5;
  assign mem[3715] = 10'd4;
  assign mem[3716] = 10'd3;
  assign mem[3717] = 10'd2;
  assign mem[3718] = 10'd3;
  assign mem[3719] = 10'd4;
  assign mem[3720] = 10'd8;
  assign mem[3721] = 10'd7;
  assign mem[3722] = 10'd6;
  assign mem[3723] = 10'd5;
  assign mem[3724] = 10'd4;
  assign mem[3725] = 10'd3;
  assign mem[3726] = 10'd2;
  assign mem[3727] = 10'd1;
  assign mem[3728] = 10'd2;
  assign mem[3729] = 10'd3;
  assign mem[3730] = 10'd7;
  assign mem[3731] = 10'd6;
  assign mem[3732] = 10'd5;
  assign mem[3733] = 10'd4;
  assign mem[3734] = 10'd3;
  assign mem[3735] = 10'd2;
  assign mem[3736] = 10'd1;
  assign mem[3737] = 10'd0;
  assign mem[3738] = 10'd1;
  assign mem[3739] = 10'd2;
  assign mem[3740] = 10'd8;
  assign mem[3741] = 10'd7;
  assign mem[3742] = 10'd6;
  assign mem[3743] = 10'd5;
  assign mem[3744] = 10'd4;
  assign mem[3745] = 10'd3;
  assign mem[3746] = 10'd2;
  assign mem[3747] = 10'd1;
  assign mem[3748] = 10'd2;
  assign mem[3749] = 10'd3;
  assign mem[3750] = 10'd9;
  assign mem[3751] = 10'd8;
  assign mem[3752] = 10'd7;
  assign mem[3753] = 10'd6;
  assign mem[3754] = 10'd5;
  assign mem[3755] = 10'd4;
  assign mem[3756] = 10'd3;
  assign mem[3757] = 10'd2;
  assign mem[3758] = 10'd3;
  assign mem[3759] = 10'd4;
  assign mem[3760] = 10'd10;
  assign mem[3761] = 10'd9;
  assign mem[3762] = 10'd8;
  assign mem[3763] = 10'd7;
  assign mem[3764] = 10'd6;
  assign mem[3765] = 10'd5;
  assign mem[3766] = 10'd4;
  assign mem[3767] = 10'd3;
  assign mem[3768] = 10'd4;
  assign mem[3769] = 10'd5;
  assign mem[3770] = 10'd11;
  assign mem[3771] = 10'd10;
  assign mem[3772] = 10'd9;
  assign mem[3773] = 10'd8;
  assign mem[3774] = 10'd7;
  assign mem[3775] = 10'd6;
  assign mem[3776] = 10'd5;
  assign mem[3777] = 10'd4;
  assign mem[3778] = 10'd5;
  assign mem[3779] = 10'd6;
  assign mem[3780] = 10'd12;
  assign mem[3781] = 10'd11;
  assign mem[3782] = 10'd10;
  assign mem[3783] = 10'd9;
  assign mem[3784] = 10'd8;
  assign mem[3785] = 10'd7;
  assign mem[3786] = 10'd6;
  assign mem[3787] = 10'd5;
  assign mem[3788] = 10'd6;
  assign mem[3789] = 10'd7;
  assign mem[3790] = 10'd13;
  assign mem[3791] = 10'd12;
  assign mem[3792] = 10'd11;
  assign mem[3793] = 10'd10;
  assign mem[3794] = 10'd9;
  assign mem[3795] = 10'd8;
  assign mem[3796] = 10'd7;
  assign mem[3797] = 10'd6;
  assign mem[3798] = 10'd7;
  assign mem[3799] = 10'd8;
  assign mem[3800] = 10'd11;
  assign mem[3801] = 10'd10;
  assign mem[3802] = 10'd9;
  assign mem[3803] = 10'd8;
  assign mem[3804] = 10'd7;
  assign mem[3805] = 10'd6;
  assign mem[3806] = 10'd5;
  assign mem[3807] = 10'd4;
  assign mem[3808] = 10'd3;
  assign mem[3809] = 10'd4;
  assign mem[3810] = 10'd10;
  assign mem[3811] = 10'd9;
  assign mem[3812] = 10'd8;
  assign mem[3813] = 10'd7;
  assign mem[3814] = 10'd6;
  assign mem[3815] = 10'd5;
  assign mem[3816] = 10'd4;
  assign mem[3817] = 10'd3;
  assign mem[3818] = 10'd2;
  assign mem[3819] = 10'd3;
  assign mem[3820] = 10'd9;
  assign mem[3821] = 10'd8;
  assign mem[3822] = 10'd7;
  assign mem[3823] = 10'd6;
  assign mem[3824] = 10'd5;
  assign mem[3825] = 10'd4;
  assign mem[3826] = 10'd3;
  assign mem[3827] = 10'd2;
  assign mem[3828] = 10'd1;
  assign mem[3829] = 10'd2;
  assign mem[3830] = 10'd8;
  assign mem[3831] = 10'd7;
  assign mem[3832] = 10'd6;
  assign mem[3833] = 10'd5;
  assign mem[3834] = 10'd4;
  assign mem[3835] = 10'd3;
  assign mem[3836] = 10'd2;
  assign mem[3837] = 10'd1;
  assign mem[3838] = 10'd0;
  assign mem[3839] = 10'd1;
  assign mem[3840] = 10'd9;
  assign mem[3841] = 10'd8;
  assign mem[3842] = 10'd7;
  assign mem[3843] = 10'd6;
  assign mem[3844] = 10'd5;
  assign mem[3845] = 10'd4;
  assign mem[3846] = 10'd3;
  assign mem[3847] = 10'd2;
  assign mem[3848] = 10'd1;
  assign mem[3849] = 10'd2;
  assign mem[3850] = 10'd10;
  assign mem[3851] = 10'd9;
  assign mem[3852] = 10'd8;
  assign mem[3853] = 10'd7;
  assign mem[3854] = 10'd6;
  assign mem[3855] = 10'd5;
  assign mem[3856] = 10'd4;
  assign mem[3857] = 10'd3;
  assign mem[3858] = 10'd2;
  assign mem[3859] = 10'd3;
  assign mem[3860] = 10'd11;
  assign mem[3861] = 10'd10;
  assign mem[3862] = 10'd9;
  assign mem[3863] = 10'd8;
  assign mem[3864] = 10'd7;
  assign mem[3865] = 10'd6;
  assign mem[3866] = 10'd5;
  assign mem[3867] = 10'd4;
  assign mem[3868] = 10'd3;
  assign mem[3869] = 10'd4;
  assign mem[3870] = 10'd12;
  assign mem[3871] = 10'd11;
  assign mem[3872] = 10'd10;
  assign mem[3873] = 10'd9;
  assign mem[3874] = 10'd8;
  assign mem[3875] = 10'd7;
  assign mem[3876] = 10'd6;
  assign mem[3877] = 10'd5;
  assign mem[3878] = 10'd4;
  assign mem[3879] = 10'd5;
  assign mem[3880] = 10'd13;
  assign mem[3881] = 10'd12;
  assign mem[3882] = 10'd11;
  assign mem[3883] = 10'd10;
  assign mem[3884] = 10'd9;
  assign mem[3885] = 10'd8;
  assign mem[3886] = 10'd7;
  assign mem[3887] = 10'd6;
  assign mem[3888] = 10'd5;
  assign mem[3889] = 10'd6;
  assign mem[3890] = 10'd14;
  assign mem[3891] = 10'd13;
  assign mem[3892] = 10'd12;
  assign mem[3893] = 10'd11;
  assign mem[3894] = 10'd10;
  assign mem[3895] = 10'd9;
  assign mem[3896] = 10'd8;
  assign mem[3897] = 10'd7;
  assign mem[3898] = 10'd6;
  assign mem[3899] = 10'd7;
  assign mem[3900] = 10'd12;
  assign mem[3901] = 10'd11;
  assign mem[3902] = 10'd10;
  assign mem[3903] = 10'd9;
  assign mem[3904] = 10'd8;
  assign mem[3905] = 10'd7;
  assign mem[3906] = 10'd6;
  assign mem[3907] = 10'd5;
  assign mem[3908] = 10'd4;
  assign mem[3909] = 10'd3;
  assign mem[3910] = 10'd11;
  assign mem[3911] = 10'd10;
  assign mem[3912] = 10'd9;
  assign mem[3913] = 10'd8;
  assign mem[3914] = 10'd7;
  assign mem[3915] = 10'd6;
  assign mem[3916] = 10'd5;
  assign mem[3917] = 10'd4;
  assign mem[3918] = 10'd3;
  assign mem[3919] = 10'd2;
  assign mem[3920] = 10'd10;
  assign mem[3921] = 10'd9;
  assign mem[3922] = 10'd8;
  assign mem[3923] = 10'd7;
  assign mem[3924] = 10'd6;
  assign mem[3925] = 10'd5;
  assign mem[3926] = 10'd4;
  assign mem[3927] = 10'd3;
  assign mem[3928] = 10'd2;
  assign mem[3929] = 10'd1;
  assign mem[3930] = 10'd9;
  assign mem[3931] = 10'd8;
  assign mem[3932] = 10'd7;
  assign mem[3933] = 10'd6;
  assign mem[3934] = 10'd5;
  assign mem[3935] = 10'd4;
  assign mem[3936] = 10'd3;
  assign mem[3937] = 10'd2;
  assign mem[3938] = 10'd1;
  assign mem[3939] = 10'd0;
  assign mem[3940] = 10'd10;
  assign mem[3941] = 10'd9;
  assign mem[3942] = 10'd8;
  assign mem[3943] = 10'd7;
  assign mem[3944] = 10'd6;
  assign mem[3945] = 10'd5;
  assign mem[3946] = 10'd4;
  assign mem[3947] = 10'd3;
  assign mem[3948] = 10'd2;
  assign mem[3949] = 10'd1;
  assign mem[3950] = 10'd11;
  assign mem[3951] = 10'd10;
  assign mem[3952] = 10'd9;
  assign mem[3953] = 10'd8;
  assign mem[3954] = 10'd7;
  assign mem[3955] = 10'd6;
  assign mem[3956] = 10'd5;
  assign mem[3957] = 10'd4;
  assign mem[3958] = 10'd3;
  assign mem[3959] = 10'd2;
  assign mem[3960] = 10'd12;
  assign mem[3961] = 10'd11;
  assign mem[3962] = 10'd10;
  assign mem[3963] = 10'd9;
  assign mem[3964] = 10'd8;
  assign mem[3965] = 10'd7;
  assign mem[3966] = 10'd6;
  assign mem[3967] = 10'd5;
  assign mem[3968] = 10'd4;
  assign mem[3969] = 10'd3;
  assign mem[3970] = 10'd13;
  assign mem[3971] = 10'd12;
  assign mem[3972] = 10'd11;
  assign mem[3973] = 10'd10;
  assign mem[3974] = 10'd9;
  assign mem[3975] = 10'd8;
  assign mem[3976] = 10'd7;
  assign mem[3977] = 10'd6;
  assign mem[3978] = 10'd5;
  assign mem[3979] = 10'd4;
  assign mem[3980] = 10'd14;
  assign mem[3981] = 10'd13;
  assign mem[3982] = 10'd12;
  assign mem[3983] = 10'd11;
  assign mem[3984] = 10'd10;
  assign mem[3985] = 10'd9;
  assign mem[3986] = 10'd8;
  assign mem[3987] = 10'd7;
  assign mem[3988] = 10'd6;
  assign mem[3989] = 10'd5;
  assign mem[3990] = 10'd15;
  assign mem[3991] = 10'd14;
  assign mem[3992] = 10'd13;
  assign mem[3993] = 10'd12;
  assign mem[3994] = 10'd11;
  assign mem[3995] = 10'd10;
  assign mem[3996] = 10'd9;
  assign mem[3997] = 10'd8;
  assign mem[3998] = 10'd7;
  assign mem[3999] = 10'd6;
  assign mem[4000] = 10'd4;
  assign mem[4001] = 10'd5;
  assign mem[4002] = 10'd6;
  assign mem[4003] = 10'd7;
  assign mem[4004] = 10'd8;
  assign mem[4005] = 10'd9;
  assign mem[4006] = 10'd10;
  assign mem[4007] = 10'd11;
  assign mem[4008] = 10'd12;
  assign mem[4009] = 10'd13;
  assign mem[4010] = 10'd3;
  assign mem[4011] = 10'd4;
  assign mem[4012] = 10'd5;
  assign mem[4013] = 10'd6;
  assign mem[4014] = 10'd7;
  assign mem[4015] = 10'd8;
  assign mem[4016] = 10'd9;
  assign mem[4017] = 10'd10;
  assign mem[4018] = 10'd11;
  assign mem[4019] = 10'd12;
  assign mem[4020] = 10'd2;
  assign mem[4021] = 10'd3;
  assign mem[4022] = 10'd4;
  assign mem[4023] = 10'd5;
  assign mem[4024] = 10'd6;
  assign mem[4025] = 10'd7;
  assign mem[4026] = 10'd8;
  assign mem[4027] = 10'd9;
  assign mem[4028] = 10'd10;
  assign mem[4029] = 10'd11;
  assign mem[4030] = 10'd1;
  assign mem[4031] = 10'd2;
  assign mem[4032] = 10'd3;
  assign mem[4033] = 10'd4;
  assign mem[4034] = 10'd5;
  assign mem[4035] = 10'd6;
  assign mem[4036] = 10'd7;
  assign mem[4037] = 10'd8;
  assign mem[4038] = 10'd9;
  assign mem[4039] = 10'd10;
  assign mem[4040] = 10'd0;
  assign mem[4041] = 10'd1;
  assign mem[4042] = 10'd2;
  assign mem[4043] = 10'd3;
  assign mem[4044] = 10'd4;
  assign mem[4045] = 10'd5;
  assign mem[4046] = 10'd6;
  assign mem[4047] = 10'd7;
  assign mem[4048] = 10'd8;
  assign mem[4049] = 10'd9;
  assign mem[4050] = 10'd1;
  assign mem[4051] = 10'd2;
  assign mem[4052] = 10'd3;
  assign mem[4053] = 10'd4;
  assign mem[4054] = 10'd5;
  assign mem[4055] = 10'd6;
  assign mem[4056] = 10'd7;
  assign mem[4057] = 10'd8;
  assign mem[4058] = 10'd9;
  assign mem[4059] = 10'd10;
  assign mem[4060] = 10'd2;
  assign mem[4061] = 10'd3;
  assign mem[4062] = 10'd4;
  assign mem[4063] = 10'd5;
  assign mem[4064] = 10'd6;
  assign mem[4065] = 10'd7;
  assign mem[4066] = 10'd8;
  assign mem[4067] = 10'd9;
  assign mem[4068] = 10'd10;
  assign mem[4069] = 10'd11;
  assign mem[4070] = 10'd3;
  assign mem[4071] = 10'd4;
  assign mem[4072] = 10'd5;
  assign mem[4073] = 10'd6;
  assign mem[4074] = 10'd7;
  assign mem[4075] = 10'd8;
  assign mem[4076] = 10'd9;
  assign mem[4077] = 10'd10;
  assign mem[4078] = 10'd11;
  assign mem[4079] = 10'd12;
  assign mem[4080] = 10'd4;
  assign mem[4081] = 10'd5;
  assign mem[4082] = 10'd6;
  assign mem[4083] = 10'd7;
  assign mem[4084] = 10'd8;
  assign mem[4085] = 10'd9;
  assign mem[4086] = 10'd10;
  assign mem[4087] = 10'd11;
  assign mem[4088] = 10'd12;
  assign mem[4089] = 10'd13;
  assign mem[4090] = 10'd5;
  assign mem[4091] = 10'd6;
  assign mem[4092] = 10'd7;
  assign mem[4093] = 10'd8;
  assign mem[4094] = 10'd9;
  assign mem[4095] = 10'd10;
  assign mem[4096] = 10'd11;
  assign mem[4097] = 10'd12;
  assign mem[4098] = 10'd13;
  assign mem[4099] = 10'd14;
  assign mem[4100] = 10'd5;
  assign mem[4101] = 10'd4;
  assign mem[4102] = 10'd5;
  assign mem[4103] = 10'd6;
  assign mem[4104] = 10'd7;
  assign mem[4105] = 10'd8;
  assign mem[4106] = 10'd9;
  assign mem[4107] = 10'd10;
  assign mem[4108] = 10'd11;
  assign mem[4109] = 10'd12;
  assign mem[4110] = 10'd4;
  assign mem[4111] = 10'd3;
  assign mem[4112] = 10'd4;
  assign mem[4113] = 10'd5;
  assign mem[4114] = 10'd6;
  assign mem[4115] = 10'd7;
  assign mem[4116] = 10'd8;
  assign mem[4117] = 10'd9;
  assign mem[4118] = 10'd10;
  assign mem[4119] = 10'd11;
  assign mem[4120] = 10'd3;
  assign mem[4121] = 10'd2;
  assign mem[4122] = 10'd3;
  assign mem[4123] = 10'd4;
  assign mem[4124] = 10'd5;
  assign mem[4125] = 10'd6;
  assign mem[4126] = 10'd7;
  assign mem[4127] = 10'd8;
  assign mem[4128] = 10'd9;
  assign mem[4129] = 10'd10;
  assign mem[4130] = 10'd2;
  assign mem[4131] = 10'd1;
  assign mem[4132] = 10'd2;
  assign mem[4133] = 10'd3;
  assign mem[4134] = 10'd4;
  assign mem[4135] = 10'd5;
  assign mem[4136] = 10'd6;
  assign mem[4137] = 10'd7;
  assign mem[4138] = 10'd8;
  assign mem[4139] = 10'd9;
  assign mem[4140] = 10'd1;
  assign mem[4141] = 10'd0;
  assign mem[4142] = 10'd1;
  assign mem[4143] = 10'd2;
  assign mem[4144] = 10'd3;
  assign mem[4145] = 10'd4;
  assign mem[4146] = 10'd5;
  assign mem[4147] = 10'd6;
  assign mem[4148] = 10'd7;
  assign mem[4149] = 10'd8;
  assign mem[4150] = 10'd2;
  assign mem[4151] = 10'd1;
  assign mem[4152] = 10'd2;
  assign mem[4153] = 10'd3;
  assign mem[4154] = 10'd4;
  assign mem[4155] = 10'd5;
  assign mem[4156] = 10'd6;
  assign mem[4157] = 10'd7;
  assign mem[4158] = 10'd8;
  assign mem[4159] = 10'd9;
  assign mem[4160] = 10'd3;
  assign mem[4161] = 10'd2;
  assign mem[4162] = 10'd3;
  assign mem[4163] = 10'd4;
  assign mem[4164] = 10'd5;
  assign mem[4165] = 10'd6;
  assign mem[4166] = 10'd7;
  assign mem[4167] = 10'd8;
  assign mem[4168] = 10'd9;
  assign mem[4169] = 10'd10;
  assign mem[4170] = 10'd4;
  assign mem[4171] = 10'd3;
  assign mem[4172] = 10'd4;
  assign mem[4173] = 10'd5;
  assign mem[4174] = 10'd6;
  assign mem[4175] = 10'd7;
  assign mem[4176] = 10'd8;
  assign mem[4177] = 10'd9;
  assign mem[4178] = 10'd10;
  assign mem[4179] = 10'd11;
  assign mem[4180] = 10'd5;
  assign mem[4181] = 10'd4;
  assign mem[4182] = 10'd5;
  assign mem[4183] = 10'd6;
  assign mem[4184] = 10'd7;
  assign mem[4185] = 10'd8;
  assign mem[4186] = 10'd9;
  assign mem[4187] = 10'd10;
  assign mem[4188] = 10'd11;
  assign mem[4189] = 10'd12;
  assign mem[4190] = 10'd6;
  assign mem[4191] = 10'd5;
  assign mem[4192] = 10'd6;
  assign mem[4193] = 10'd7;
  assign mem[4194] = 10'd8;
  assign mem[4195] = 10'd9;
  assign mem[4196] = 10'd10;
  assign mem[4197] = 10'd11;
  assign mem[4198] = 10'd12;
  assign mem[4199] = 10'd13;
  assign mem[4200] = 10'd6;
  assign mem[4201] = 10'd5;
  assign mem[4202] = 10'd4;
  assign mem[4203] = 10'd5;
  assign mem[4204] = 10'd6;
  assign mem[4205] = 10'd7;
  assign mem[4206] = 10'd8;
  assign mem[4207] = 10'd9;
  assign mem[4208] = 10'd10;
  assign mem[4209] = 10'd11;
  assign mem[4210] = 10'd5;
  assign mem[4211] = 10'd4;
  assign mem[4212] = 10'd3;
  assign mem[4213] = 10'd4;
  assign mem[4214] = 10'd5;
  assign mem[4215] = 10'd6;
  assign mem[4216] = 10'd7;
  assign mem[4217] = 10'd8;
  assign mem[4218] = 10'd9;
  assign mem[4219] = 10'd10;
  assign mem[4220] = 10'd4;
  assign mem[4221] = 10'd3;
  assign mem[4222] = 10'd2;
  assign mem[4223] = 10'd3;
  assign mem[4224] = 10'd4;
  assign mem[4225] = 10'd5;
  assign mem[4226] = 10'd6;
  assign mem[4227] = 10'd7;
  assign mem[4228] = 10'd8;
  assign mem[4229] = 10'd9;
  assign mem[4230] = 10'd3;
  assign mem[4231] = 10'd2;
  assign mem[4232] = 10'd1;
  assign mem[4233] = 10'd2;
  assign mem[4234] = 10'd3;
  assign mem[4235] = 10'd4;
  assign mem[4236] = 10'd5;
  assign mem[4237] = 10'd6;
  assign mem[4238] = 10'd7;
  assign mem[4239] = 10'd8;
  assign mem[4240] = 10'd2;
  assign mem[4241] = 10'd1;
  assign mem[4242] = 10'd0;
  assign mem[4243] = 10'd1;
  assign mem[4244] = 10'd2;
  assign mem[4245] = 10'd3;
  assign mem[4246] = 10'd4;
  assign mem[4247] = 10'd5;
  assign mem[4248] = 10'd6;
  assign mem[4249] = 10'd7;
  assign mem[4250] = 10'd3;
  assign mem[4251] = 10'd2;
  assign mem[4252] = 10'd1;
  assign mem[4253] = 10'd2;
  assign mem[4254] = 10'd3;
  assign mem[4255] = 10'd4;
  assign mem[4256] = 10'd5;
  assign mem[4257] = 10'd6;
  assign mem[4258] = 10'd7;
  assign mem[4259] = 10'd8;
  assign mem[4260] = 10'd4;
  assign mem[4261] = 10'd3;
  assign mem[4262] = 10'd2;
  assign mem[4263] = 10'd3;
  assign mem[4264] = 10'd4;
  assign mem[4265] = 10'd5;
  assign mem[4266] = 10'd6;
  assign mem[4267] = 10'd7;
  assign mem[4268] = 10'd8;
  assign mem[4269] = 10'd9;
  assign mem[4270] = 10'd5;
  assign mem[4271] = 10'd4;
  assign mem[4272] = 10'd3;
  assign mem[4273] = 10'd4;
  assign mem[4274] = 10'd5;
  assign mem[4275] = 10'd6;
  assign mem[4276] = 10'd7;
  assign mem[4277] = 10'd8;
  assign mem[4278] = 10'd9;
  assign mem[4279] = 10'd10;
  assign mem[4280] = 10'd6;
  assign mem[4281] = 10'd5;
  assign mem[4282] = 10'd4;
  assign mem[4283] = 10'd5;
  assign mem[4284] = 10'd6;
  assign mem[4285] = 10'd7;
  assign mem[4286] = 10'd8;
  assign mem[4287] = 10'd9;
  assign mem[4288] = 10'd10;
  assign mem[4289] = 10'd11;
  assign mem[4290] = 10'd7;
  assign mem[4291] = 10'd6;
  assign mem[4292] = 10'd5;
  assign mem[4293] = 10'd6;
  assign mem[4294] = 10'd7;
  assign mem[4295] = 10'd8;
  assign mem[4296] = 10'd9;
  assign mem[4297] = 10'd10;
  assign mem[4298] = 10'd11;
  assign mem[4299] = 10'd12;
  assign mem[4300] = 10'd7;
  assign mem[4301] = 10'd6;
  assign mem[4302] = 10'd5;
  assign mem[4303] = 10'd4;
  assign mem[4304] = 10'd5;
  assign mem[4305] = 10'd6;
  assign mem[4306] = 10'd7;
  assign mem[4307] = 10'd8;
  assign mem[4308] = 10'd9;
  assign mem[4309] = 10'd10;
  assign mem[4310] = 10'd6;
  assign mem[4311] = 10'd5;
  assign mem[4312] = 10'd4;
  assign mem[4313] = 10'd3;
  assign mem[4314] = 10'd4;
  assign mem[4315] = 10'd5;
  assign mem[4316] = 10'd6;
  assign mem[4317] = 10'd7;
  assign mem[4318] = 10'd8;
  assign mem[4319] = 10'd9;
  assign mem[4320] = 10'd5;
  assign mem[4321] = 10'd4;
  assign mem[4322] = 10'd3;
  assign mem[4323] = 10'd2;
  assign mem[4324] = 10'd3;
  assign mem[4325] = 10'd4;
  assign mem[4326] = 10'd5;
  assign mem[4327] = 10'd6;
  assign mem[4328] = 10'd7;
  assign mem[4329] = 10'd8;
  assign mem[4330] = 10'd4;
  assign mem[4331] = 10'd3;
  assign mem[4332] = 10'd2;
  assign mem[4333] = 10'd1;
  assign mem[4334] = 10'd2;
  assign mem[4335] = 10'd3;
  assign mem[4336] = 10'd4;
  assign mem[4337] = 10'd5;
  assign mem[4338] = 10'd6;
  assign mem[4339] = 10'd7;
  assign mem[4340] = 10'd3;
  assign mem[4341] = 10'd2;
  assign mem[4342] = 10'd1;
  assign mem[4343] = 10'd0;
  assign mem[4344] = 10'd1;
  assign mem[4345] = 10'd2;
  assign mem[4346] = 10'd3;
  assign mem[4347] = 10'd4;
  assign mem[4348] = 10'd5;
  assign mem[4349] = 10'd6;
  assign mem[4350] = 10'd4;
  assign mem[4351] = 10'd3;
  assign mem[4352] = 10'd2;
  assign mem[4353] = 10'd1;
  assign mem[4354] = 10'd2;
  assign mem[4355] = 10'd3;
  assign mem[4356] = 10'd4;
  assign mem[4357] = 10'd5;
  assign mem[4358] = 10'd6;
  assign mem[4359] = 10'd7;
  assign mem[4360] = 10'd5;
  assign mem[4361] = 10'd4;
  assign mem[4362] = 10'd3;
  assign mem[4363] = 10'd2;
  assign mem[4364] = 10'd3;
  assign mem[4365] = 10'd4;
  assign mem[4366] = 10'd5;
  assign mem[4367] = 10'd6;
  assign mem[4368] = 10'd7;
  assign mem[4369] = 10'd8;
  assign mem[4370] = 10'd6;
  assign mem[4371] = 10'd5;
  assign mem[4372] = 10'd4;
  assign mem[4373] = 10'd3;
  assign mem[4374] = 10'd4;
  assign mem[4375] = 10'd5;
  assign mem[4376] = 10'd6;
  assign mem[4377] = 10'd7;
  assign mem[4378] = 10'd8;
  assign mem[4379] = 10'd9;
  assign mem[4380] = 10'd7;
  assign mem[4381] = 10'd6;
  assign mem[4382] = 10'd5;
  assign mem[4383] = 10'd4;
  assign mem[4384] = 10'd5;
  assign mem[4385] = 10'd6;
  assign mem[4386] = 10'd7;
  assign mem[4387] = 10'd8;
  assign mem[4388] = 10'd9;
  assign mem[4389] = 10'd10;
  assign mem[4390] = 10'd8;
  assign mem[4391] = 10'd7;
  assign mem[4392] = 10'd6;
  assign mem[4393] = 10'd5;
  assign mem[4394] = 10'd6;
  assign mem[4395] = 10'd7;
  assign mem[4396] = 10'd8;
  assign mem[4397] = 10'd9;
  assign mem[4398] = 10'd10;
  assign mem[4399] = 10'd11;
  assign mem[4400] = 10'd8;
  assign mem[4401] = 10'd7;
  assign mem[4402] = 10'd6;
  assign mem[4403] = 10'd5;
  assign mem[4404] = 10'd4;
  assign mem[4405] = 10'd5;
  assign mem[4406] = 10'd6;
  assign mem[4407] = 10'd7;
  assign mem[4408] = 10'd8;
  assign mem[4409] = 10'd9;
  assign mem[4410] = 10'd7;
  assign mem[4411] = 10'd6;
  assign mem[4412] = 10'd5;
  assign mem[4413] = 10'd4;
  assign mem[4414] = 10'd3;
  assign mem[4415] = 10'd4;
  assign mem[4416] = 10'd5;
  assign mem[4417] = 10'd6;
  assign mem[4418] = 10'd7;
  assign mem[4419] = 10'd8;
  assign mem[4420] = 10'd6;
  assign mem[4421] = 10'd5;
  assign mem[4422] = 10'd4;
  assign mem[4423] = 10'd3;
  assign mem[4424] = 10'd2;
  assign mem[4425] = 10'd3;
  assign mem[4426] = 10'd4;
  assign mem[4427] = 10'd5;
  assign mem[4428] = 10'd6;
  assign mem[4429] = 10'd7;
  assign mem[4430] = 10'd5;
  assign mem[4431] = 10'd4;
  assign mem[4432] = 10'd3;
  assign mem[4433] = 10'd2;
  assign mem[4434] = 10'd1;
  assign mem[4435] = 10'd2;
  assign mem[4436] = 10'd3;
  assign mem[4437] = 10'd4;
  assign mem[4438] = 10'd5;
  assign mem[4439] = 10'd6;
  assign mem[4440] = 10'd4;
  assign mem[4441] = 10'd3;
  assign mem[4442] = 10'd2;
  assign mem[4443] = 10'd1;
  assign mem[4444] = 10'd0;
  assign mem[4445] = 10'd1;
  assign mem[4446] = 10'd2;
  assign mem[4447] = 10'd3;
  assign mem[4448] = 10'd4;
  assign mem[4449] = 10'd5;
  assign mem[4450] = 10'd5;
  assign mem[4451] = 10'd4;
  assign mem[4452] = 10'd3;
  assign mem[4453] = 10'd2;
  assign mem[4454] = 10'd1;
  assign mem[4455] = 10'd2;
  assign mem[4456] = 10'd3;
  assign mem[4457] = 10'd4;
  assign mem[4458] = 10'd5;
  assign mem[4459] = 10'd6;
  assign mem[4460] = 10'd6;
  assign mem[4461] = 10'd5;
  assign mem[4462] = 10'd4;
  assign mem[4463] = 10'd3;
  assign mem[4464] = 10'd2;
  assign mem[4465] = 10'd3;
  assign mem[4466] = 10'd4;
  assign mem[4467] = 10'd5;
  assign mem[4468] = 10'd6;
  assign mem[4469] = 10'd7;
  assign mem[4470] = 10'd7;
  assign mem[4471] = 10'd6;
  assign mem[4472] = 10'd5;
  assign mem[4473] = 10'd4;
  assign mem[4474] = 10'd3;
  assign mem[4475] = 10'd4;
  assign mem[4476] = 10'd5;
  assign mem[4477] = 10'd6;
  assign mem[4478] = 10'd7;
  assign mem[4479] = 10'd8;
  assign mem[4480] = 10'd8;
  assign mem[4481] = 10'd7;
  assign mem[4482] = 10'd6;
  assign mem[4483] = 10'd5;
  assign mem[4484] = 10'd4;
  assign mem[4485] = 10'd5;
  assign mem[4486] = 10'd6;
  assign mem[4487] = 10'd7;
  assign mem[4488] = 10'd8;
  assign mem[4489] = 10'd9;
  assign mem[4490] = 10'd9;
  assign mem[4491] = 10'd8;
  assign mem[4492] = 10'd7;
  assign mem[4493] = 10'd6;
  assign mem[4494] = 10'd5;
  assign mem[4495] = 10'd6;
  assign mem[4496] = 10'd7;
  assign mem[4497] = 10'd8;
  assign mem[4498] = 10'd9;
  assign mem[4499] = 10'd10;
  assign mem[4500] = 10'd9;
  assign mem[4501] = 10'd8;
  assign mem[4502] = 10'd7;
  assign mem[4503] = 10'd6;
  assign mem[4504] = 10'd5;
  assign mem[4505] = 10'd4;
  assign mem[4506] = 10'd5;
  assign mem[4507] = 10'd6;
  assign mem[4508] = 10'd7;
  assign mem[4509] = 10'd8;
  assign mem[4510] = 10'd8;
  assign mem[4511] = 10'd7;
  assign mem[4512] = 10'd6;
  assign mem[4513] = 10'd5;
  assign mem[4514] = 10'd4;
  assign mem[4515] = 10'd3;
  assign mem[4516] = 10'd4;
  assign mem[4517] = 10'd5;
  assign mem[4518] = 10'd6;
  assign mem[4519] = 10'd7;
  assign mem[4520] = 10'd7;
  assign mem[4521] = 10'd6;
  assign mem[4522] = 10'd5;
  assign mem[4523] = 10'd4;
  assign mem[4524] = 10'd3;
  assign mem[4525] = 10'd2;
  assign mem[4526] = 10'd3;
  assign mem[4527] = 10'd4;
  assign mem[4528] = 10'd5;
  assign mem[4529] = 10'd6;
  assign mem[4530] = 10'd6;
  assign mem[4531] = 10'd5;
  assign mem[4532] = 10'd4;
  assign mem[4533] = 10'd3;
  assign mem[4534] = 10'd2;
  assign mem[4535] = 10'd1;
  assign mem[4536] = 10'd2;
  assign mem[4537] = 10'd3;
  assign mem[4538] = 10'd4;
  assign mem[4539] = 10'd5;
  assign mem[4540] = 10'd5;
  assign mem[4541] = 10'd4;
  assign mem[4542] = 10'd3;
  assign mem[4543] = 10'd2;
  assign mem[4544] = 10'd1;
  assign mem[4545] = 10'd0;
  assign mem[4546] = 10'd1;
  assign mem[4547] = 10'd2;
  assign mem[4548] = 10'd3;
  assign mem[4549] = 10'd4;
  assign mem[4550] = 10'd6;
  assign mem[4551] = 10'd5;
  assign mem[4552] = 10'd4;
  assign mem[4553] = 10'd3;
  assign mem[4554] = 10'd2;
  assign mem[4555] = 10'd1;
  assign mem[4556] = 10'd2;
  assign mem[4557] = 10'd3;
  assign mem[4558] = 10'd4;
  assign mem[4559] = 10'd5;
  assign mem[4560] = 10'd7;
  assign mem[4561] = 10'd6;
  assign mem[4562] = 10'd5;
  assign mem[4563] = 10'd4;
  assign mem[4564] = 10'd3;
  assign mem[4565] = 10'd2;
  assign mem[4566] = 10'd3;
  assign mem[4567] = 10'd4;
  assign mem[4568] = 10'd5;
  assign mem[4569] = 10'd6;
  assign mem[4570] = 10'd8;
  assign mem[4571] = 10'd7;
  assign mem[4572] = 10'd6;
  assign mem[4573] = 10'd5;
  assign mem[4574] = 10'd4;
  assign mem[4575] = 10'd3;
  assign mem[4576] = 10'd4;
  assign mem[4577] = 10'd5;
  assign mem[4578] = 10'd6;
  assign mem[4579] = 10'd7;
  assign mem[4580] = 10'd9;
  assign mem[4581] = 10'd8;
  assign mem[4582] = 10'd7;
  assign mem[4583] = 10'd6;
  assign mem[4584] = 10'd5;
  assign mem[4585] = 10'd4;
  assign mem[4586] = 10'd5;
  assign mem[4587] = 10'd6;
  assign mem[4588] = 10'd7;
  assign mem[4589] = 10'd8;
  assign mem[4590] = 10'd10;
  assign mem[4591] = 10'd9;
  assign mem[4592] = 10'd8;
  assign mem[4593] = 10'd7;
  assign mem[4594] = 10'd6;
  assign mem[4595] = 10'd5;
  assign mem[4596] = 10'd6;
  assign mem[4597] = 10'd7;
  assign mem[4598] = 10'd8;
  assign mem[4599] = 10'd9;
  assign mem[4600] = 10'd10;
  assign mem[4601] = 10'd9;
  assign mem[4602] = 10'd8;
  assign mem[4603] = 10'd7;
  assign mem[4604] = 10'd6;
  assign mem[4605] = 10'd5;
  assign mem[4606] = 10'd4;
  assign mem[4607] = 10'd5;
  assign mem[4608] = 10'd6;
  assign mem[4609] = 10'd7;
  assign mem[4610] = 10'd9;
  assign mem[4611] = 10'd8;
  assign mem[4612] = 10'd7;
  assign mem[4613] = 10'd6;
  assign mem[4614] = 10'd5;
  assign mem[4615] = 10'd4;
  assign mem[4616] = 10'd3;
  assign mem[4617] = 10'd4;
  assign mem[4618] = 10'd5;
  assign mem[4619] = 10'd6;
  assign mem[4620] = 10'd8;
  assign mem[4621] = 10'd7;
  assign mem[4622] = 10'd6;
  assign mem[4623] = 10'd5;
  assign mem[4624] = 10'd4;
  assign mem[4625] = 10'd3;
  assign mem[4626] = 10'd2;
  assign mem[4627] = 10'd3;
  assign mem[4628] = 10'd4;
  assign mem[4629] = 10'd5;
  assign mem[4630] = 10'd7;
  assign mem[4631] = 10'd6;
  assign mem[4632] = 10'd5;
  assign mem[4633] = 10'd4;
  assign mem[4634] = 10'd3;
  assign mem[4635] = 10'd2;
  assign mem[4636] = 10'd1;
  assign mem[4637] = 10'd2;
  assign mem[4638] = 10'd3;
  assign mem[4639] = 10'd4;
  assign mem[4640] = 10'd6;
  assign mem[4641] = 10'd5;
  assign mem[4642] = 10'd4;
  assign mem[4643] = 10'd3;
  assign mem[4644] = 10'd2;
  assign mem[4645] = 10'd1;
  assign mem[4646] = 10'd0;
  assign mem[4647] = 10'd1;
  assign mem[4648] = 10'd2;
  assign mem[4649] = 10'd3;
  assign mem[4650] = 10'd7;
  assign mem[4651] = 10'd6;
  assign mem[4652] = 10'd5;
  assign mem[4653] = 10'd4;
  assign mem[4654] = 10'd3;
  assign mem[4655] = 10'd2;
  assign mem[4656] = 10'd1;
  assign mem[4657] = 10'd2;
  assign mem[4658] = 10'd3;
  assign mem[4659] = 10'd4;
  assign mem[4660] = 10'd8;
  assign mem[4661] = 10'd7;
  assign mem[4662] = 10'd6;
  assign mem[4663] = 10'd5;
  assign mem[4664] = 10'd4;
  assign mem[4665] = 10'd3;
  assign mem[4666] = 10'd2;
  assign mem[4667] = 10'd3;
  assign mem[4668] = 10'd4;
  assign mem[4669] = 10'd5;
  assign mem[4670] = 10'd9;
  assign mem[4671] = 10'd8;
  assign mem[4672] = 10'd7;
  assign mem[4673] = 10'd6;
  assign mem[4674] = 10'd5;
  assign mem[4675] = 10'd4;
  assign mem[4676] = 10'd3;
  assign mem[4677] = 10'd4;
  assign mem[4678] = 10'd5;
  assign mem[4679] = 10'd6;
  assign mem[4680] = 10'd10;
  assign mem[4681] = 10'd9;
  assign mem[4682] = 10'd8;
  assign mem[4683] = 10'd7;
  assign mem[4684] = 10'd6;
  assign mem[4685] = 10'd5;
  assign mem[4686] = 10'd4;
  assign mem[4687] = 10'd5;
  assign mem[4688] = 10'd6;
  assign mem[4689] = 10'd7;
  assign mem[4690] = 10'd11;
  assign mem[4691] = 10'd10;
  assign mem[4692] = 10'd9;
  assign mem[4693] = 10'd8;
  assign mem[4694] = 10'd7;
  assign mem[4695] = 10'd6;
  assign mem[4696] = 10'd5;
  assign mem[4697] = 10'd6;
  assign mem[4698] = 10'd7;
  assign mem[4699] = 10'd8;
  assign mem[4700] = 10'd11;
  assign mem[4701] = 10'd10;
  assign mem[4702] = 10'd9;
  assign mem[4703] = 10'd8;
  assign mem[4704] = 10'd7;
  assign mem[4705] = 10'd6;
  assign mem[4706] = 10'd5;
  assign mem[4707] = 10'd4;
  assign mem[4708] = 10'd5;
  assign mem[4709] = 10'd6;
  assign mem[4710] = 10'd10;
  assign mem[4711] = 10'd9;
  assign mem[4712] = 10'd8;
  assign mem[4713] = 10'd7;
  assign mem[4714] = 10'd6;
  assign mem[4715] = 10'd5;
  assign mem[4716] = 10'd4;
  assign mem[4717] = 10'd3;
  assign mem[4718] = 10'd4;
  assign mem[4719] = 10'd5;
  assign mem[4720] = 10'd9;
  assign mem[4721] = 10'd8;
  assign mem[4722] = 10'd7;
  assign mem[4723] = 10'd6;
  assign mem[4724] = 10'd5;
  assign mem[4725] = 10'd4;
  assign mem[4726] = 10'd3;
  assign mem[4727] = 10'd2;
  assign mem[4728] = 10'd3;
  assign mem[4729] = 10'd4;
  assign mem[4730] = 10'd8;
  assign mem[4731] = 10'd7;
  assign mem[4732] = 10'd6;
  assign mem[4733] = 10'd5;
  assign mem[4734] = 10'd4;
  assign mem[4735] = 10'd3;
  assign mem[4736] = 10'd2;
  assign mem[4737] = 10'd1;
  assign mem[4738] = 10'd2;
  assign mem[4739] = 10'd3;
  assign mem[4740] = 10'd7;
  assign mem[4741] = 10'd6;
  assign mem[4742] = 10'd5;
  assign mem[4743] = 10'd4;
  assign mem[4744] = 10'd3;
  assign mem[4745] = 10'd2;
  assign mem[4746] = 10'd1;
  assign mem[4747] = 10'd0;
  assign mem[4748] = 10'd1;
  assign mem[4749] = 10'd2;
  assign mem[4750] = 10'd8;
  assign mem[4751] = 10'd7;
  assign mem[4752] = 10'd6;
  assign mem[4753] = 10'd5;
  assign mem[4754] = 10'd4;
  assign mem[4755] = 10'd3;
  assign mem[4756] = 10'd2;
  assign mem[4757] = 10'd1;
  assign mem[4758] = 10'd2;
  assign mem[4759] = 10'd3;
  assign mem[4760] = 10'd9;
  assign mem[4761] = 10'd8;
  assign mem[4762] = 10'd7;
  assign mem[4763] = 10'd6;
  assign mem[4764] = 10'd5;
  assign mem[4765] = 10'd4;
  assign mem[4766] = 10'd3;
  assign mem[4767] = 10'd2;
  assign mem[4768] = 10'd3;
  assign mem[4769] = 10'd4;
  assign mem[4770] = 10'd10;
  assign mem[4771] = 10'd9;
  assign mem[4772] = 10'd8;
  assign mem[4773] = 10'd7;
  assign mem[4774] = 10'd6;
  assign mem[4775] = 10'd5;
  assign mem[4776] = 10'd4;
  assign mem[4777] = 10'd3;
  assign mem[4778] = 10'd4;
  assign mem[4779] = 10'd5;
  assign mem[4780] = 10'd11;
  assign mem[4781] = 10'd10;
  assign mem[4782] = 10'd9;
  assign mem[4783] = 10'd8;
  assign mem[4784] = 10'd7;
  assign mem[4785] = 10'd6;
  assign mem[4786] = 10'd5;
  assign mem[4787] = 10'd4;
  assign mem[4788] = 10'd5;
  assign mem[4789] = 10'd6;
  assign mem[4790] = 10'd12;
  assign mem[4791] = 10'd11;
  assign mem[4792] = 10'd10;
  assign mem[4793] = 10'd9;
  assign mem[4794] = 10'd8;
  assign mem[4795] = 10'd7;
  assign mem[4796] = 10'd6;
  assign mem[4797] = 10'd5;
  assign mem[4798] = 10'd6;
  assign mem[4799] = 10'd7;
  assign mem[4800] = 10'd12;
  assign mem[4801] = 10'd11;
  assign mem[4802] = 10'd10;
  assign mem[4803] = 10'd9;
  assign mem[4804] = 10'd8;
  assign mem[4805] = 10'd7;
  assign mem[4806] = 10'd6;
  assign mem[4807] = 10'd5;
  assign mem[4808] = 10'd4;
  assign mem[4809] = 10'd5;
  assign mem[4810] = 10'd11;
  assign mem[4811] = 10'd10;
  assign mem[4812] = 10'd9;
  assign mem[4813] = 10'd8;
  assign mem[4814] = 10'd7;
  assign mem[4815] = 10'd6;
  assign mem[4816] = 10'd5;
  assign mem[4817] = 10'd4;
  assign mem[4818] = 10'd3;
  assign mem[4819] = 10'd4;
  assign mem[4820] = 10'd10;
  assign mem[4821] = 10'd9;
  assign mem[4822] = 10'd8;
  assign mem[4823] = 10'd7;
  assign mem[4824] = 10'd6;
  assign mem[4825] = 10'd5;
  assign mem[4826] = 10'd4;
  assign mem[4827] = 10'd3;
  assign mem[4828] = 10'd2;
  assign mem[4829] = 10'd3;
  assign mem[4830] = 10'd9;
  assign mem[4831] = 10'd8;
  assign mem[4832] = 10'd7;
  assign mem[4833] = 10'd6;
  assign mem[4834] = 10'd5;
  assign mem[4835] = 10'd4;
  assign mem[4836] = 10'd3;
  assign mem[4837] = 10'd2;
  assign mem[4838] = 10'd1;
  assign mem[4839] = 10'd2;
  assign mem[4840] = 10'd8;
  assign mem[4841] = 10'd7;
  assign mem[4842] = 10'd6;
  assign mem[4843] = 10'd5;
  assign mem[4844] = 10'd4;
  assign mem[4845] = 10'd3;
  assign mem[4846] = 10'd2;
  assign mem[4847] = 10'd1;
  assign mem[4848] = 10'd0;
  assign mem[4849] = 10'd1;
  assign mem[4850] = 10'd9;
  assign mem[4851] = 10'd8;
  assign mem[4852] = 10'd7;
  assign mem[4853] = 10'd6;
  assign mem[4854] = 10'd5;
  assign mem[4855] = 10'd4;
  assign mem[4856] = 10'd3;
  assign mem[4857] = 10'd2;
  assign mem[4858] = 10'd1;
  assign mem[4859] = 10'd2;
  assign mem[4860] = 10'd10;
  assign mem[4861] = 10'd9;
  assign mem[4862] = 10'd8;
  assign mem[4863] = 10'd7;
  assign mem[4864] = 10'd6;
  assign mem[4865] = 10'd5;
  assign mem[4866] = 10'd4;
  assign mem[4867] = 10'd3;
  assign mem[4868] = 10'd2;
  assign mem[4869] = 10'd3;
  assign mem[4870] = 10'd11;
  assign mem[4871] = 10'd10;
  assign mem[4872] = 10'd9;
  assign mem[4873] = 10'd8;
  assign mem[4874] = 10'd7;
  assign mem[4875] = 10'd6;
  assign mem[4876] = 10'd5;
  assign mem[4877] = 10'd4;
  assign mem[4878] = 10'd3;
  assign mem[4879] = 10'd4;
  assign mem[4880] = 10'd12;
  assign mem[4881] = 10'd11;
  assign mem[4882] = 10'd10;
  assign mem[4883] = 10'd9;
  assign mem[4884] = 10'd8;
  assign mem[4885] = 10'd7;
  assign mem[4886] = 10'd6;
  assign mem[4887] = 10'd5;
  assign mem[4888] = 10'd4;
  assign mem[4889] = 10'd5;
  assign mem[4890] = 10'd13;
  assign mem[4891] = 10'd12;
  assign mem[4892] = 10'd11;
  assign mem[4893] = 10'd10;
  assign mem[4894] = 10'd9;
  assign mem[4895] = 10'd8;
  assign mem[4896] = 10'd7;
  assign mem[4897] = 10'd6;
  assign mem[4898] = 10'd5;
  assign mem[4899] = 10'd6;
  assign mem[4900] = 10'd13;
  assign mem[4901] = 10'd12;
  assign mem[4902] = 10'd11;
  assign mem[4903] = 10'd10;
  assign mem[4904] = 10'd9;
  assign mem[4905] = 10'd8;
  assign mem[4906] = 10'd7;
  assign mem[4907] = 10'd6;
  assign mem[4908] = 10'd5;
  assign mem[4909] = 10'd4;
  assign mem[4910] = 10'd12;
  assign mem[4911] = 10'd11;
  assign mem[4912] = 10'd10;
  assign mem[4913] = 10'd9;
  assign mem[4914] = 10'd8;
  assign mem[4915] = 10'd7;
  assign mem[4916] = 10'd6;
  assign mem[4917] = 10'd5;
  assign mem[4918] = 10'd4;
  assign mem[4919] = 10'd3;
  assign mem[4920] = 10'd11;
  assign mem[4921] = 10'd10;
  assign mem[4922] = 10'd9;
  assign mem[4923] = 10'd8;
  assign mem[4924] = 10'd7;
  assign mem[4925] = 10'd6;
  assign mem[4926] = 10'd5;
  assign mem[4927] = 10'd4;
  assign mem[4928] = 10'd3;
  assign mem[4929] = 10'd2;
  assign mem[4930] = 10'd10;
  assign mem[4931] = 10'd9;
  assign mem[4932] = 10'd8;
  assign mem[4933] = 10'd7;
  assign mem[4934] = 10'd6;
  assign mem[4935] = 10'd5;
  assign mem[4936] = 10'd4;
  assign mem[4937] = 10'd3;
  assign mem[4938] = 10'd2;
  assign mem[4939] = 10'd1;
  assign mem[4940] = 10'd9;
  assign mem[4941] = 10'd8;
  assign mem[4942] = 10'd7;
  assign mem[4943] = 10'd6;
  assign mem[4944] = 10'd5;
  assign mem[4945] = 10'd4;
  assign mem[4946] = 10'd3;
  assign mem[4947] = 10'd2;
  assign mem[4948] = 10'd1;
  assign mem[4949] = 10'd0;
  assign mem[4950] = 10'd10;
  assign mem[4951] = 10'd9;
  assign mem[4952] = 10'd8;
  assign mem[4953] = 10'd7;
  assign mem[4954] = 10'd6;
  assign mem[4955] = 10'd5;
  assign mem[4956] = 10'd4;
  assign mem[4957] = 10'd3;
  assign mem[4958] = 10'd2;
  assign mem[4959] = 10'd1;
  assign mem[4960] = 10'd11;
  assign mem[4961] = 10'd10;
  assign mem[4962] = 10'd9;
  assign mem[4963] = 10'd8;
  assign mem[4964] = 10'd7;
  assign mem[4965] = 10'd6;
  assign mem[4966] = 10'd5;
  assign mem[4967] = 10'd4;
  assign mem[4968] = 10'd3;
  assign mem[4969] = 10'd2;
  assign mem[4970] = 10'd12;
  assign mem[4971] = 10'd11;
  assign mem[4972] = 10'd10;
  assign mem[4973] = 10'd9;
  assign mem[4974] = 10'd8;
  assign mem[4975] = 10'd7;
  assign mem[4976] = 10'd6;
  assign mem[4977] = 10'd5;
  assign mem[4978] = 10'd4;
  assign mem[4979] = 10'd3;
  assign mem[4980] = 10'd13;
  assign mem[4981] = 10'd12;
  assign mem[4982] = 10'd11;
  assign mem[4983] = 10'd10;
  assign mem[4984] = 10'd9;
  assign mem[4985] = 10'd8;
  assign mem[4986] = 10'd7;
  assign mem[4987] = 10'd6;
  assign mem[4988] = 10'd5;
  assign mem[4989] = 10'd4;
  assign mem[4990] = 10'd14;
  assign mem[4991] = 10'd13;
  assign mem[4992] = 10'd12;
  assign mem[4993] = 10'd11;
  assign mem[4994] = 10'd10;
  assign mem[4995] = 10'd9;
  assign mem[4996] = 10'd8;
  assign mem[4997] = 10'd7;
  assign mem[4998] = 10'd6;
  assign mem[4999] = 10'd5;
  assign mem[5000] = 10'd5;
  assign mem[5001] = 10'd6;
  assign mem[5002] = 10'd7;
  assign mem[5003] = 10'd8;
  assign mem[5004] = 10'd9;
  assign mem[5005] = 10'd10;
  assign mem[5006] = 10'd11;
  assign mem[5007] = 10'd12;
  assign mem[5008] = 10'd13;
  assign mem[5009] = 10'd14;
  assign mem[5010] = 10'd4;
  assign mem[5011] = 10'd5;
  assign mem[5012] = 10'd6;
  assign mem[5013] = 10'd7;
  assign mem[5014] = 10'd8;
  assign mem[5015] = 10'd9;
  assign mem[5016] = 10'd10;
  assign mem[5017] = 10'd11;
  assign mem[5018] = 10'd12;
  assign mem[5019] = 10'd13;
  assign mem[5020] = 10'd3;
  assign mem[5021] = 10'd4;
  assign mem[5022] = 10'd5;
  assign mem[5023] = 10'd6;
  assign mem[5024] = 10'd7;
  assign mem[5025] = 10'd8;
  assign mem[5026] = 10'd9;
  assign mem[5027] = 10'd10;
  assign mem[5028] = 10'd11;
  assign mem[5029] = 10'd12;
  assign mem[5030] = 10'd2;
  assign mem[5031] = 10'd3;
  assign mem[5032] = 10'd4;
  assign mem[5033] = 10'd5;
  assign mem[5034] = 10'd6;
  assign mem[5035] = 10'd7;
  assign mem[5036] = 10'd8;
  assign mem[5037] = 10'd9;
  assign mem[5038] = 10'd10;
  assign mem[5039] = 10'd11;
  assign mem[5040] = 10'd1;
  assign mem[5041] = 10'd2;
  assign mem[5042] = 10'd3;
  assign mem[5043] = 10'd4;
  assign mem[5044] = 10'd5;
  assign mem[5045] = 10'd6;
  assign mem[5046] = 10'd7;
  assign mem[5047] = 10'd8;
  assign mem[5048] = 10'd9;
  assign mem[5049] = 10'd10;
  assign mem[5050] = 10'd0;
  assign mem[5051] = 10'd1;
  assign mem[5052] = 10'd2;
  assign mem[5053] = 10'd3;
  assign mem[5054] = 10'd4;
  assign mem[5055] = 10'd5;
  assign mem[5056] = 10'd6;
  assign mem[5057] = 10'd7;
  assign mem[5058] = 10'd8;
  assign mem[5059] = 10'd9;
  assign mem[5060] = 10'd1;
  assign mem[5061] = 10'd2;
  assign mem[5062] = 10'd3;
  assign mem[5063] = 10'd4;
  assign mem[5064] = 10'd5;
  assign mem[5065] = 10'd6;
  assign mem[5066] = 10'd7;
  assign mem[5067] = 10'd8;
  assign mem[5068] = 10'd9;
  assign mem[5069] = 10'd10;
  assign mem[5070] = 10'd2;
  assign mem[5071] = 10'd3;
  assign mem[5072] = 10'd4;
  assign mem[5073] = 10'd5;
  assign mem[5074] = 10'd6;
  assign mem[5075] = 10'd7;
  assign mem[5076] = 10'd8;
  assign mem[5077] = 10'd9;
  assign mem[5078] = 10'd10;
  assign mem[5079] = 10'd11;
  assign mem[5080] = 10'd3;
  assign mem[5081] = 10'd4;
  assign mem[5082] = 10'd5;
  assign mem[5083] = 10'd6;
  assign mem[5084] = 10'd7;
  assign mem[5085] = 10'd8;
  assign mem[5086] = 10'd9;
  assign mem[5087] = 10'd10;
  assign mem[5088] = 10'd11;
  assign mem[5089] = 10'd12;
  assign mem[5090] = 10'd4;
  assign mem[5091] = 10'd5;
  assign mem[5092] = 10'd6;
  assign mem[5093] = 10'd7;
  assign mem[5094] = 10'd8;
  assign mem[5095] = 10'd9;
  assign mem[5096] = 10'd10;
  assign mem[5097] = 10'd11;
  assign mem[5098] = 10'd12;
  assign mem[5099] = 10'd13;
  assign mem[5100] = 10'd6;
  assign mem[5101] = 10'd5;
  assign mem[5102] = 10'd6;
  assign mem[5103] = 10'd7;
  assign mem[5104] = 10'd8;
  assign mem[5105] = 10'd9;
  assign mem[5106] = 10'd10;
  assign mem[5107] = 10'd11;
  assign mem[5108] = 10'd12;
  assign mem[5109] = 10'd13;
  assign mem[5110] = 10'd5;
  assign mem[5111] = 10'd4;
  assign mem[5112] = 10'd5;
  assign mem[5113] = 10'd6;
  assign mem[5114] = 10'd7;
  assign mem[5115] = 10'd8;
  assign mem[5116] = 10'd9;
  assign mem[5117] = 10'd10;
  assign mem[5118] = 10'd11;
  assign mem[5119] = 10'd12;
  assign mem[5120] = 10'd4;
  assign mem[5121] = 10'd3;
  assign mem[5122] = 10'd4;
  assign mem[5123] = 10'd5;
  assign mem[5124] = 10'd6;
  assign mem[5125] = 10'd7;
  assign mem[5126] = 10'd8;
  assign mem[5127] = 10'd9;
  assign mem[5128] = 10'd10;
  assign mem[5129] = 10'd11;
  assign mem[5130] = 10'd3;
  assign mem[5131] = 10'd2;
  assign mem[5132] = 10'd3;
  assign mem[5133] = 10'd4;
  assign mem[5134] = 10'd5;
  assign mem[5135] = 10'd6;
  assign mem[5136] = 10'd7;
  assign mem[5137] = 10'd8;
  assign mem[5138] = 10'd9;
  assign mem[5139] = 10'd10;
  assign mem[5140] = 10'd2;
  assign mem[5141] = 10'd1;
  assign mem[5142] = 10'd2;
  assign mem[5143] = 10'd3;
  assign mem[5144] = 10'd4;
  assign mem[5145] = 10'd5;
  assign mem[5146] = 10'd6;
  assign mem[5147] = 10'd7;
  assign mem[5148] = 10'd8;
  assign mem[5149] = 10'd9;
  assign mem[5150] = 10'd1;
  assign mem[5151] = 10'd0;
  assign mem[5152] = 10'd1;
  assign mem[5153] = 10'd2;
  assign mem[5154] = 10'd3;
  assign mem[5155] = 10'd4;
  assign mem[5156] = 10'd5;
  assign mem[5157] = 10'd6;
  assign mem[5158] = 10'd7;
  assign mem[5159] = 10'd8;
  assign mem[5160] = 10'd2;
  assign mem[5161] = 10'd1;
  assign mem[5162] = 10'd2;
  assign mem[5163] = 10'd3;
  assign mem[5164] = 10'd4;
  assign mem[5165] = 10'd5;
  assign mem[5166] = 10'd6;
  assign mem[5167] = 10'd7;
  assign mem[5168] = 10'd8;
  assign mem[5169] = 10'd9;
  assign mem[5170] = 10'd3;
  assign mem[5171] = 10'd2;
  assign mem[5172] = 10'd3;
  assign mem[5173] = 10'd4;
  assign mem[5174] = 10'd5;
  assign mem[5175] = 10'd6;
  assign mem[5176] = 10'd7;
  assign mem[5177] = 10'd8;
  assign mem[5178] = 10'd9;
  assign mem[5179] = 10'd10;
  assign mem[5180] = 10'd4;
  assign mem[5181] = 10'd3;
  assign mem[5182] = 10'd4;
  assign mem[5183] = 10'd5;
  assign mem[5184] = 10'd6;
  assign mem[5185] = 10'd7;
  assign mem[5186] = 10'd8;
  assign mem[5187] = 10'd9;
  assign mem[5188] = 10'd10;
  assign mem[5189] = 10'd11;
  assign mem[5190] = 10'd5;
  assign mem[5191] = 10'd4;
  assign mem[5192] = 10'd5;
  assign mem[5193] = 10'd6;
  assign mem[5194] = 10'd7;
  assign mem[5195] = 10'd8;
  assign mem[5196] = 10'd9;
  assign mem[5197] = 10'd10;
  assign mem[5198] = 10'd11;
  assign mem[5199] = 10'd12;
  assign mem[5200] = 10'd7;
  assign mem[5201] = 10'd6;
  assign mem[5202] = 10'd5;
  assign mem[5203] = 10'd6;
  assign mem[5204] = 10'd7;
  assign mem[5205] = 10'd8;
  assign mem[5206] = 10'd9;
  assign mem[5207] = 10'd10;
  assign mem[5208] = 10'd11;
  assign mem[5209] = 10'd12;
  assign mem[5210] = 10'd6;
  assign mem[5211] = 10'd5;
  assign mem[5212] = 10'd4;
  assign mem[5213] = 10'd5;
  assign mem[5214] = 10'd6;
  assign mem[5215] = 10'd7;
  assign mem[5216] = 10'd8;
  assign mem[5217] = 10'd9;
  assign mem[5218] = 10'd10;
  assign mem[5219] = 10'd11;
  assign mem[5220] = 10'd5;
  assign mem[5221] = 10'd4;
  assign mem[5222] = 10'd3;
  assign mem[5223] = 10'd4;
  assign mem[5224] = 10'd5;
  assign mem[5225] = 10'd6;
  assign mem[5226] = 10'd7;
  assign mem[5227] = 10'd8;
  assign mem[5228] = 10'd9;
  assign mem[5229] = 10'd10;
  assign mem[5230] = 10'd4;
  assign mem[5231] = 10'd3;
  assign mem[5232] = 10'd2;
  assign mem[5233] = 10'd3;
  assign mem[5234] = 10'd4;
  assign mem[5235] = 10'd5;
  assign mem[5236] = 10'd6;
  assign mem[5237] = 10'd7;
  assign mem[5238] = 10'd8;
  assign mem[5239] = 10'd9;
  assign mem[5240] = 10'd3;
  assign mem[5241] = 10'd2;
  assign mem[5242] = 10'd1;
  assign mem[5243] = 10'd2;
  assign mem[5244] = 10'd3;
  assign mem[5245] = 10'd4;
  assign mem[5246] = 10'd5;
  assign mem[5247] = 10'd6;
  assign mem[5248] = 10'd7;
  assign mem[5249] = 10'd8;
  assign mem[5250] = 10'd2;
  assign mem[5251] = 10'd1;
  assign mem[5252] = 10'd0;
  assign mem[5253] = 10'd1;
  assign mem[5254] = 10'd2;
  assign mem[5255] = 10'd3;
  assign mem[5256] = 10'd4;
  assign mem[5257] = 10'd5;
  assign mem[5258] = 10'd6;
  assign mem[5259] = 10'd7;
  assign mem[5260] = 10'd3;
  assign mem[5261] = 10'd2;
  assign mem[5262] = 10'd1;
  assign mem[5263] = 10'd2;
  assign mem[5264] = 10'd3;
  assign mem[5265] = 10'd4;
  assign mem[5266] = 10'd5;
  assign mem[5267] = 10'd6;
  assign mem[5268] = 10'd7;
  assign mem[5269] = 10'd8;
  assign mem[5270] = 10'd4;
  assign mem[5271] = 10'd3;
  assign mem[5272] = 10'd2;
  assign mem[5273] = 10'd3;
  assign mem[5274] = 10'd4;
  assign mem[5275] = 10'd5;
  assign mem[5276] = 10'd6;
  assign mem[5277] = 10'd7;
  assign mem[5278] = 10'd8;
  assign mem[5279] = 10'd9;
  assign mem[5280] = 10'd5;
  assign mem[5281] = 10'd4;
  assign mem[5282] = 10'd3;
  assign mem[5283] = 10'd4;
  assign mem[5284] = 10'd5;
  assign mem[5285] = 10'd6;
  assign mem[5286] = 10'd7;
  assign mem[5287] = 10'd8;
  assign mem[5288] = 10'd9;
  assign mem[5289] = 10'd10;
  assign mem[5290] = 10'd6;
  assign mem[5291] = 10'd5;
  assign mem[5292] = 10'd4;
  assign mem[5293] = 10'd5;
  assign mem[5294] = 10'd6;
  assign mem[5295] = 10'd7;
  assign mem[5296] = 10'd8;
  assign mem[5297] = 10'd9;
  assign mem[5298] = 10'd10;
  assign mem[5299] = 10'd11;
  assign mem[5300] = 10'd8;
  assign mem[5301] = 10'd7;
  assign mem[5302] = 10'd6;
  assign mem[5303] = 10'd5;
  assign mem[5304] = 10'd6;
  assign mem[5305] = 10'd7;
  assign mem[5306] = 10'd8;
  assign mem[5307] = 10'd9;
  assign mem[5308] = 10'd10;
  assign mem[5309] = 10'd11;
  assign mem[5310] = 10'd7;
  assign mem[5311] = 10'd6;
  assign mem[5312] = 10'd5;
  assign mem[5313] = 10'd4;
  assign mem[5314] = 10'd5;
  assign mem[5315] = 10'd6;
  assign mem[5316] = 10'd7;
  assign mem[5317] = 10'd8;
  assign mem[5318] = 10'd9;
  assign mem[5319] = 10'd10;
  assign mem[5320] = 10'd6;
  assign mem[5321] = 10'd5;
  assign mem[5322] = 10'd4;
  assign mem[5323] = 10'd3;
  assign mem[5324] = 10'd4;
  assign mem[5325] = 10'd5;
  assign mem[5326] = 10'd6;
  assign mem[5327] = 10'd7;
  assign mem[5328] = 10'd8;
  assign mem[5329] = 10'd9;
  assign mem[5330] = 10'd5;
  assign mem[5331] = 10'd4;
  assign mem[5332] = 10'd3;
  assign mem[5333] = 10'd2;
  assign mem[5334] = 10'd3;
  assign mem[5335] = 10'd4;
  assign mem[5336] = 10'd5;
  assign mem[5337] = 10'd6;
  assign mem[5338] = 10'd7;
  assign mem[5339] = 10'd8;
  assign mem[5340] = 10'd4;
  assign mem[5341] = 10'd3;
  assign mem[5342] = 10'd2;
  assign mem[5343] = 10'd1;
  assign mem[5344] = 10'd2;
  assign mem[5345] = 10'd3;
  assign mem[5346] = 10'd4;
  assign mem[5347] = 10'd5;
  assign mem[5348] = 10'd6;
  assign mem[5349] = 10'd7;
  assign mem[5350] = 10'd3;
  assign mem[5351] = 10'd2;
  assign mem[5352] = 10'd1;
  assign mem[5353] = 10'd0;
  assign mem[5354] = 10'd1;
  assign mem[5355] = 10'd2;
  assign mem[5356] = 10'd3;
  assign mem[5357] = 10'd4;
  assign mem[5358] = 10'd5;
  assign mem[5359] = 10'd6;
  assign mem[5360] = 10'd4;
  assign mem[5361] = 10'd3;
  assign mem[5362] = 10'd2;
  assign mem[5363] = 10'd1;
  assign mem[5364] = 10'd2;
  assign mem[5365] = 10'd3;
  assign mem[5366] = 10'd4;
  assign mem[5367] = 10'd5;
  assign mem[5368] = 10'd6;
  assign mem[5369] = 10'd7;
  assign mem[5370] = 10'd5;
  assign mem[5371] = 10'd4;
  assign mem[5372] = 10'd3;
  assign mem[5373] = 10'd2;
  assign mem[5374] = 10'd3;
  assign mem[5375] = 10'd4;
  assign mem[5376] = 10'd5;
  assign mem[5377] = 10'd6;
  assign mem[5378] = 10'd7;
  assign mem[5379] = 10'd8;
  assign mem[5380] = 10'd6;
  assign mem[5381] = 10'd5;
  assign mem[5382] = 10'd4;
  assign mem[5383] = 10'd3;
  assign mem[5384] = 10'd4;
  assign mem[5385] = 10'd5;
  assign mem[5386] = 10'd6;
  assign mem[5387] = 10'd7;
  assign mem[5388] = 10'd8;
  assign mem[5389] = 10'd9;
  assign mem[5390] = 10'd7;
  assign mem[5391] = 10'd6;
  assign mem[5392] = 10'd5;
  assign mem[5393] = 10'd4;
  assign mem[5394] = 10'd5;
  assign mem[5395] = 10'd6;
  assign mem[5396] = 10'd7;
  assign mem[5397] = 10'd8;
  assign mem[5398] = 10'd9;
  assign mem[5399] = 10'd10;
  assign mem[5400] = 10'd9;
  assign mem[5401] = 10'd8;
  assign mem[5402] = 10'd7;
  assign mem[5403] = 10'd6;
  assign mem[5404] = 10'd5;
  assign mem[5405] = 10'd6;
  assign mem[5406] = 10'd7;
  assign mem[5407] = 10'd8;
  assign mem[5408] = 10'd9;
  assign mem[5409] = 10'd10;
  assign mem[5410] = 10'd8;
  assign mem[5411] = 10'd7;
  assign mem[5412] = 10'd6;
  assign mem[5413] = 10'd5;
  assign mem[5414] = 10'd4;
  assign mem[5415] = 10'd5;
  assign mem[5416] = 10'd6;
  assign mem[5417] = 10'd7;
  assign mem[5418] = 10'd8;
  assign mem[5419] = 10'd9;
  assign mem[5420] = 10'd7;
  assign mem[5421] = 10'd6;
  assign mem[5422] = 10'd5;
  assign mem[5423] = 10'd4;
  assign mem[5424] = 10'd3;
  assign mem[5425] = 10'd4;
  assign mem[5426] = 10'd5;
  assign mem[5427] = 10'd6;
  assign mem[5428] = 10'd7;
  assign mem[5429] = 10'd8;
  assign mem[5430] = 10'd6;
  assign mem[5431] = 10'd5;
  assign mem[5432] = 10'd4;
  assign mem[5433] = 10'd3;
  assign mem[5434] = 10'd2;
  assign mem[5435] = 10'd3;
  assign mem[5436] = 10'd4;
  assign mem[5437] = 10'd5;
  assign mem[5438] = 10'd6;
  assign mem[5439] = 10'd7;
  assign mem[5440] = 10'd5;
  assign mem[5441] = 10'd4;
  assign mem[5442] = 10'd3;
  assign mem[5443] = 10'd2;
  assign mem[5444] = 10'd1;
  assign mem[5445] = 10'd2;
  assign mem[5446] = 10'd3;
  assign mem[5447] = 10'd4;
  assign mem[5448] = 10'd5;
  assign mem[5449] = 10'd6;
  assign mem[5450] = 10'd4;
  assign mem[5451] = 10'd3;
  assign mem[5452] = 10'd2;
  assign mem[5453] = 10'd1;
  assign mem[5454] = 10'd0;
  assign mem[5455] = 10'd1;
  assign mem[5456] = 10'd2;
  assign mem[5457] = 10'd3;
  assign mem[5458] = 10'd4;
  assign mem[5459] = 10'd5;
  assign mem[5460] = 10'd5;
  assign mem[5461] = 10'd4;
  assign mem[5462] = 10'd3;
  assign mem[5463] = 10'd2;
  assign mem[5464] = 10'd1;
  assign mem[5465] = 10'd2;
  assign mem[5466] = 10'd3;
  assign mem[5467] = 10'd4;
  assign mem[5468] = 10'd5;
  assign mem[5469] = 10'd6;
  assign mem[5470] = 10'd6;
  assign mem[5471] = 10'd5;
  assign mem[5472] = 10'd4;
  assign mem[5473] = 10'd3;
  assign mem[5474] = 10'd2;
  assign mem[5475] = 10'd3;
  assign mem[5476] = 10'd4;
  assign mem[5477] = 10'd5;
  assign mem[5478] = 10'd6;
  assign mem[5479] = 10'd7;
  assign mem[5480] = 10'd7;
  assign mem[5481] = 10'd6;
  assign mem[5482] = 10'd5;
  assign mem[5483] = 10'd4;
  assign mem[5484] = 10'd3;
  assign mem[5485] = 10'd4;
  assign mem[5486] = 10'd5;
  assign mem[5487] = 10'd6;
  assign mem[5488] = 10'd7;
  assign mem[5489] = 10'd8;
  assign mem[5490] = 10'd8;
  assign mem[5491] = 10'd7;
  assign mem[5492] = 10'd6;
  assign mem[5493] = 10'd5;
  assign mem[5494] = 10'd4;
  assign mem[5495] = 10'd5;
  assign mem[5496] = 10'd6;
  assign mem[5497] = 10'd7;
  assign mem[5498] = 10'd8;
  assign mem[5499] = 10'd9;
  assign mem[5500] = 10'd10;
  assign mem[5501] = 10'd9;
  assign mem[5502] = 10'd8;
  assign mem[5503] = 10'd7;
  assign mem[5504] = 10'd6;
  assign mem[5505] = 10'd5;
  assign mem[5506] = 10'd6;
  assign mem[5507] = 10'd7;
  assign mem[5508] = 10'd8;
  assign mem[5509] = 10'd9;
  assign mem[5510] = 10'd9;
  assign mem[5511] = 10'd8;
  assign mem[5512] = 10'd7;
  assign mem[5513] = 10'd6;
  assign mem[5514] = 10'd5;
  assign mem[5515] = 10'd4;
  assign mem[5516] = 10'd5;
  assign mem[5517] = 10'd6;
  assign mem[5518] = 10'd7;
  assign mem[5519] = 10'd8;
  assign mem[5520] = 10'd8;
  assign mem[5521] = 10'd7;
  assign mem[5522] = 10'd6;
  assign mem[5523] = 10'd5;
  assign mem[5524] = 10'd4;
  assign mem[5525] = 10'd3;
  assign mem[5526] = 10'd4;
  assign mem[5527] = 10'd5;
  assign mem[5528] = 10'd6;
  assign mem[5529] = 10'd7;
  assign mem[5530] = 10'd7;
  assign mem[5531] = 10'd6;
  assign mem[5532] = 10'd5;
  assign mem[5533] = 10'd4;
  assign mem[5534] = 10'd3;
  assign mem[5535] = 10'd2;
  assign mem[5536] = 10'd3;
  assign mem[5537] = 10'd4;
  assign mem[5538] = 10'd5;
  assign mem[5539] = 10'd6;
  assign mem[5540] = 10'd6;
  assign mem[5541] = 10'd5;
  assign mem[5542] = 10'd4;
  assign mem[5543] = 10'd3;
  assign mem[5544] = 10'd2;
  assign mem[5545] = 10'd1;
  assign mem[5546] = 10'd2;
  assign mem[5547] = 10'd3;
  assign mem[5548] = 10'd4;
  assign mem[5549] = 10'd5;
  assign mem[5550] = 10'd5;
  assign mem[5551] = 10'd4;
  assign mem[5552] = 10'd3;
  assign mem[5553] = 10'd2;
  assign mem[5554] = 10'd1;
  assign mem[5555] = 10'd0;
  assign mem[5556] = 10'd1;
  assign mem[5557] = 10'd2;
  assign mem[5558] = 10'd3;
  assign mem[5559] = 10'd4;
  assign mem[5560] = 10'd6;
  assign mem[5561] = 10'd5;
  assign mem[5562] = 10'd4;
  assign mem[5563] = 10'd3;
  assign mem[5564] = 10'd2;
  assign mem[5565] = 10'd1;
  assign mem[5566] = 10'd2;
  assign mem[5567] = 10'd3;
  assign mem[5568] = 10'd4;
  assign mem[5569] = 10'd5;
  assign mem[5570] = 10'd7;
  assign mem[5571] = 10'd6;
  assign mem[5572] = 10'd5;
  assign mem[5573] = 10'd4;
  assign mem[5574] = 10'd3;
  assign mem[5575] = 10'd2;
  assign mem[5576] = 10'd3;
  assign mem[5577] = 10'd4;
  assign mem[5578] = 10'd5;
  assign mem[5579] = 10'd6;
  assign mem[5580] = 10'd8;
  assign mem[5581] = 10'd7;
  assign mem[5582] = 10'd6;
  assign mem[5583] = 10'd5;
  assign mem[5584] = 10'd4;
  assign mem[5585] = 10'd3;
  assign mem[5586] = 10'd4;
  assign mem[5587] = 10'd5;
  assign mem[5588] = 10'd6;
  assign mem[5589] = 10'd7;
  assign mem[5590] = 10'd9;
  assign mem[5591] = 10'd8;
  assign mem[5592] = 10'd7;
  assign mem[5593] = 10'd6;
  assign mem[5594] = 10'd5;
  assign mem[5595] = 10'd4;
  assign mem[5596] = 10'd5;
  assign mem[5597] = 10'd6;
  assign mem[5598] = 10'd7;
  assign mem[5599] = 10'd8;
  assign mem[5600] = 10'd11;
  assign mem[5601] = 10'd10;
  assign mem[5602] = 10'd9;
  assign mem[5603] = 10'd8;
  assign mem[5604] = 10'd7;
  assign mem[5605] = 10'd6;
  assign mem[5606] = 10'd5;
  assign mem[5607] = 10'd6;
  assign mem[5608] = 10'd7;
  assign mem[5609] = 10'd8;
  assign mem[5610] = 10'd10;
  assign mem[5611] = 10'd9;
  assign mem[5612] = 10'd8;
  assign mem[5613] = 10'd7;
  assign mem[5614] = 10'd6;
  assign mem[5615] = 10'd5;
  assign mem[5616] = 10'd4;
  assign mem[5617] = 10'd5;
  assign mem[5618] = 10'd6;
  assign mem[5619] = 10'd7;
  assign mem[5620] = 10'd9;
  assign mem[5621] = 10'd8;
  assign mem[5622] = 10'd7;
  assign mem[5623] = 10'd6;
  assign mem[5624] = 10'd5;
  assign mem[5625] = 10'd4;
  assign mem[5626] = 10'd3;
  assign mem[5627] = 10'd4;
  assign mem[5628] = 10'd5;
  assign mem[5629] = 10'd6;
  assign mem[5630] = 10'd8;
  assign mem[5631] = 10'd7;
  assign mem[5632] = 10'd6;
  assign mem[5633] = 10'd5;
  assign mem[5634] = 10'd4;
  assign mem[5635] = 10'd3;
  assign mem[5636] = 10'd2;
  assign mem[5637] = 10'd3;
  assign mem[5638] = 10'd4;
  assign mem[5639] = 10'd5;
  assign mem[5640] = 10'd7;
  assign mem[5641] = 10'd6;
  assign mem[5642] = 10'd5;
  assign mem[5643] = 10'd4;
  assign mem[5644] = 10'd3;
  assign mem[5645] = 10'd2;
  assign mem[5646] = 10'd1;
  assign mem[5647] = 10'd2;
  assign mem[5648] = 10'd3;
  assign mem[5649] = 10'd4;
  assign mem[5650] = 10'd6;
  assign mem[5651] = 10'd5;
  assign mem[5652] = 10'd4;
  assign mem[5653] = 10'd3;
  assign mem[5654] = 10'd2;
  assign mem[5655] = 10'd1;
  assign mem[5656] = 10'd0;
  assign mem[5657] = 10'd1;
  assign mem[5658] = 10'd2;
  assign mem[5659] = 10'd3;
  assign mem[5660] = 10'd7;
  assign mem[5661] = 10'd6;
  assign mem[5662] = 10'd5;
  assign mem[5663] = 10'd4;
  assign mem[5664] = 10'd3;
  assign mem[5665] = 10'd2;
  assign mem[5666] = 10'd1;
  assign mem[5667] = 10'd2;
  assign mem[5668] = 10'd3;
  assign mem[5669] = 10'd4;
  assign mem[5670] = 10'd8;
  assign mem[5671] = 10'd7;
  assign mem[5672] = 10'd6;
  assign mem[5673] = 10'd5;
  assign mem[5674] = 10'd4;
  assign mem[5675] = 10'd3;
  assign mem[5676] = 10'd2;
  assign mem[5677] = 10'd3;
  assign mem[5678] = 10'd4;
  assign mem[5679] = 10'd5;
  assign mem[5680] = 10'd9;
  assign mem[5681] = 10'd8;
  assign mem[5682] = 10'd7;
  assign mem[5683] = 10'd6;
  assign mem[5684] = 10'd5;
  assign mem[5685] = 10'd4;
  assign mem[5686] = 10'd3;
  assign mem[5687] = 10'd4;
  assign mem[5688] = 10'd5;
  assign mem[5689] = 10'd6;
  assign mem[5690] = 10'd10;
  assign mem[5691] = 10'd9;
  assign mem[5692] = 10'd8;
  assign mem[5693] = 10'd7;
  assign mem[5694] = 10'd6;
  assign mem[5695] = 10'd5;
  assign mem[5696] = 10'd4;
  assign mem[5697] = 10'd5;
  assign mem[5698] = 10'd6;
  assign mem[5699] = 10'd7;
  assign mem[5700] = 10'd12;
  assign mem[5701] = 10'd11;
  assign mem[5702] = 10'd10;
  assign mem[5703] = 10'd9;
  assign mem[5704] = 10'd8;
  assign mem[5705] = 10'd7;
  assign mem[5706] = 10'd6;
  assign mem[5707] = 10'd5;
  assign mem[5708] = 10'd6;
  assign mem[5709] = 10'd7;
  assign mem[5710] = 10'd11;
  assign mem[5711] = 10'd10;
  assign mem[5712] = 10'd9;
  assign mem[5713] = 10'd8;
  assign mem[5714] = 10'd7;
  assign mem[5715] = 10'd6;
  assign mem[5716] = 10'd5;
  assign mem[5717] = 10'd4;
  assign mem[5718] = 10'd5;
  assign mem[5719] = 10'd6;
  assign mem[5720] = 10'd10;
  assign mem[5721] = 10'd9;
  assign mem[5722] = 10'd8;
  assign mem[5723] = 10'd7;
  assign mem[5724] = 10'd6;
  assign mem[5725] = 10'd5;
  assign mem[5726] = 10'd4;
  assign mem[5727] = 10'd3;
  assign mem[5728] = 10'd4;
  assign mem[5729] = 10'd5;
  assign mem[5730] = 10'd9;
  assign mem[5731] = 10'd8;
  assign mem[5732] = 10'd7;
  assign mem[5733] = 10'd6;
  assign mem[5734] = 10'd5;
  assign mem[5735] = 10'd4;
  assign mem[5736] = 10'd3;
  assign mem[5737] = 10'd2;
  assign mem[5738] = 10'd3;
  assign mem[5739] = 10'd4;
  assign mem[5740] = 10'd8;
  assign mem[5741] = 10'd7;
  assign mem[5742] = 10'd6;
  assign mem[5743] = 10'd5;
  assign mem[5744] = 10'd4;
  assign mem[5745] = 10'd3;
  assign mem[5746] = 10'd2;
  assign mem[5747] = 10'd1;
  assign mem[5748] = 10'd2;
  assign mem[5749] = 10'd3;
  assign mem[5750] = 10'd7;
  assign mem[5751] = 10'd6;
  assign mem[5752] = 10'd5;
  assign mem[5753] = 10'd4;
  assign mem[5754] = 10'd3;
  assign mem[5755] = 10'd2;
  assign mem[5756] = 10'd1;
  assign mem[5757] = 10'd0;
  assign mem[5758] = 10'd1;
  assign mem[5759] = 10'd2;
  assign mem[5760] = 10'd8;
  assign mem[5761] = 10'd7;
  assign mem[5762] = 10'd6;
  assign mem[5763] = 10'd5;
  assign mem[5764] = 10'd4;
  assign mem[5765] = 10'd3;
  assign mem[5766] = 10'd2;
  assign mem[5767] = 10'd1;
  assign mem[5768] = 10'd2;
  assign mem[5769] = 10'd3;
  assign mem[5770] = 10'd9;
  assign mem[5771] = 10'd8;
  assign mem[5772] = 10'd7;
  assign mem[5773] = 10'd6;
  assign mem[5774] = 10'd5;
  assign mem[5775] = 10'd4;
  assign mem[5776] = 10'd3;
  assign mem[5777] = 10'd2;
  assign mem[5778] = 10'd3;
  assign mem[5779] = 10'd4;
  assign mem[5780] = 10'd10;
  assign mem[5781] = 10'd9;
  assign mem[5782] = 10'd8;
  assign mem[5783] = 10'd7;
  assign mem[5784] = 10'd6;
  assign mem[5785] = 10'd5;
  assign mem[5786] = 10'd4;
  assign mem[5787] = 10'd3;
  assign mem[5788] = 10'd4;
  assign mem[5789] = 10'd5;
  assign mem[5790] = 10'd11;
  assign mem[5791] = 10'd10;
  assign mem[5792] = 10'd9;
  assign mem[5793] = 10'd8;
  assign mem[5794] = 10'd7;
  assign mem[5795] = 10'd6;
  assign mem[5796] = 10'd5;
  assign mem[5797] = 10'd4;
  assign mem[5798] = 10'd5;
  assign mem[5799] = 10'd6;
  assign mem[5800] = 10'd13;
  assign mem[5801] = 10'd12;
  assign mem[5802] = 10'd11;
  assign mem[5803] = 10'd10;
  assign mem[5804] = 10'd9;
  assign mem[5805] = 10'd8;
  assign mem[5806] = 10'd7;
  assign mem[5807] = 10'd6;
  assign mem[5808] = 10'd5;
  assign mem[5809] = 10'd6;
  assign mem[5810] = 10'd12;
  assign mem[5811] = 10'd11;
  assign mem[5812] = 10'd10;
  assign mem[5813] = 10'd9;
  assign mem[5814] = 10'd8;
  assign mem[5815] = 10'd7;
  assign mem[5816] = 10'd6;
  assign mem[5817] = 10'd5;
  assign mem[5818] = 10'd4;
  assign mem[5819] = 10'd5;
  assign mem[5820] = 10'd11;
  assign mem[5821] = 10'd10;
  assign mem[5822] = 10'd9;
  assign mem[5823] = 10'd8;
  assign mem[5824] = 10'd7;
  assign mem[5825] = 10'd6;
  assign mem[5826] = 10'd5;
  assign mem[5827] = 10'd4;
  assign mem[5828] = 10'd3;
  assign mem[5829] = 10'd4;
  assign mem[5830] = 10'd10;
  assign mem[5831] = 10'd9;
  assign mem[5832] = 10'd8;
  assign mem[5833] = 10'd7;
  assign mem[5834] = 10'd6;
  assign mem[5835] = 10'd5;
  assign mem[5836] = 10'd4;
  assign mem[5837] = 10'd3;
  assign mem[5838] = 10'd2;
  assign mem[5839] = 10'd3;
  assign mem[5840] = 10'd9;
  assign mem[5841] = 10'd8;
  assign mem[5842] = 10'd7;
  assign mem[5843] = 10'd6;
  assign mem[5844] = 10'd5;
  assign mem[5845] = 10'd4;
  assign mem[5846] = 10'd3;
  assign mem[5847] = 10'd2;
  assign mem[5848] = 10'd1;
  assign mem[5849] = 10'd2;
  assign mem[5850] = 10'd8;
  assign mem[5851] = 10'd7;
  assign mem[5852] = 10'd6;
  assign mem[5853] = 10'd5;
  assign mem[5854] = 10'd4;
  assign mem[5855] = 10'd3;
  assign mem[5856] = 10'd2;
  assign mem[5857] = 10'd1;
  assign mem[5858] = 10'd0;
  assign mem[5859] = 10'd1;
  assign mem[5860] = 10'd9;
  assign mem[5861] = 10'd8;
  assign mem[5862] = 10'd7;
  assign mem[5863] = 10'd6;
  assign mem[5864] = 10'd5;
  assign mem[5865] = 10'd4;
  assign mem[5866] = 10'd3;
  assign mem[5867] = 10'd2;
  assign mem[5868] = 10'd1;
  assign mem[5869] = 10'd2;
  assign mem[5870] = 10'd10;
  assign mem[5871] = 10'd9;
  assign mem[5872] = 10'd8;
  assign mem[5873] = 10'd7;
  assign mem[5874] = 10'd6;
  assign mem[5875] = 10'd5;
  assign mem[5876] = 10'd4;
  assign mem[5877] = 10'd3;
  assign mem[5878] = 10'd2;
  assign mem[5879] = 10'd3;
  assign mem[5880] = 10'd11;
  assign mem[5881] = 10'd10;
  assign mem[5882] = 10'd9;
  assign mem[5883] = 10'd8;
  assign mem[5884] = 10'd7;
  assign mem[5885] = 10'd6;
  assign mem[5886] = 10'd5;
  assign mem[5887] = 10'd4;
  assign mem[5888] = 10'd3;
  assign mem[5889] = 10'd4;
  assign mem[5890] = 10'd12;
  assign mem[5891] = 10'd11;
  assign mem[5892] = 10'd10;
  assign mem[5893] = 10'd9;
  assign mem[5894] = 10'd8;
  assign mem[5895] = 10'd7;
  assign mem[5896] = 10'd6;
  assign mem[5897] = 10'd5;
  assign mem[5898] = 10'd4;
  assign mem[5899] = 10'd5;
  assign mem[5900] = 10'd14;
  assign mem[5901] = 10'd13;
  assign mem[5902] = 10'd12;
  assign mem[5903] = 10'd11;
  assign mem[5904] = 10'd10;
  assign mem[5905] = 10'd9;
  assign mem[5906] = 10'd8;
  assign mem[5907] = 10'd7;
  assign mem[5908] = 10'd6;
  assign mem[5909] = 10'd5;
  assign mem[5910] = 10'd13;
  assign mem[5911] = 10'd12;
  assign mem[5912] = 10'd11;
  assign mem[5913] = 10'd10;
  assign mem[5914] = 10'd9;
  assign mem[5915] = 10'd8;
  assign mem[5916] = 10'd7;
  assign mem[5917] = 10'd6;
  assign mem[5918] = 10'd5;
  assign mem[5919] = 10'd4;
  assign mem[5920] = 10'd12;
  assign mem[5921] = 10'd11;
  assign mem[5922] = 10'd10;
  assign mem[5923] = 10'd9;
  assign mem[5924] = 10'd8;
  assign mem[5925] = 10'd7;
  assign mem[5926] = 10'd6;
  assign mem[5927] = 10'd5;
  assign mem[5928] = 10'd4;
  assign mem[5929] = 10'd3;
  assign mem[5930] = 10'd11;
  assign mem[5931] = 10'd10;
  assign mem[5932] = 10'd9;
  assign mem[5933] = 10'd8;
  assign mem[5934] = 10'd7;
  assign mem[5935] = 10'd6;
  assign mem[5936] = 10'd5;
  assign mem[5937] = 10'd4;
  assign mem[5938] = 10'd3;
  assign mem[5939] = 10'd2;
  assign mem[5940] = 10'd10;
  assign mem[5941] = 10'd9;
  assign mem[5942] = 10'd8;
  assign mem[5943] = 10'd7;
  assign mem[5944] = 10'd6;
  assign mem[5945] = 10'd5;
  assign mem[5946] = 10'd4;
  assign mem[5947] = 10'd3;
  assign mem[5948] = 10'd2;
  assign mem[5949] = 10'd1;
  assign mem[5950] = 10'd9;
  assign mem[5951] = 10'd8;
  assign mem[5952] = 10'd7;
  assign mem[5953] = 10'd6;
  assign mem[5954] = 10'd5;
  assign mem[5955] = 10'd4;
  assign mem[5956] = 10'd3;
  assign mem[5957] = 10'd2;
  assign mem[5958] = 10'd1;
  assign mem[5959] = 10'd0;
  assign mem[5960] = 10'd10;
  assign mem[5961] = 10'd9;
  assign mem[5962] = 10'd8;
  assign mem[5963] = 10'd7;
  assign mem[5964] = 10'd6;
  assign mem[5965] = 10'd5;
  assign mem[5966] = 10'd4;
  assign mem[5967] = 10'd3;
  assign mem[5968] = 10'd2;
  assign mem[5969] = 10'd1;
  assign mem[5970] = 10'd11;
  assign mem[5971] = 10'd10;
  assign mem[5972] = 10'd9;
  assign mem[5973] = 10'd8;
  assign mem[5974] = 10'd7;
  assign mem[5975] = 10'd6;
  assign mem[5976] = 10'd5;
  assign mem[5977] = 10'd4;
  assign mem[5978] = 10'd3;
  assign mem[5979] = 10'd2;
  assign mem[5980] = 10'd12;
  assign mem[5981] = 10'd11;
  assign mem[5982] = 10'd10;
  assign mem[5983] = 10'd9;
  assign mem[5984] = 10'd8;
  assign mem[5985] = 10'd7;
  assign mem[5986] = 10'd6;
  assign mem[5987] = 10'd5;
  assign mem[5988] = 10'd4;
  assign mem[5989] = 10'd3;
  assign mem[5990] = 10'd13;
  assign mem[5991] = 10'd12;
  assign mem[5992] = 10'd11;
  assign mem[5993] = 10'd10;
  assign mem[5994] = 10'd9;
  assign mem[5995] = 10'd8;
  assign mem[5996] = 10'd7;
  assign mem[5997] = 10'd6;
  assign mem[5998] = 10'd5;
  assign mem[5999] = 10'd4;
  assign mem[6000] = 10'd6;
  assign mem[6001] = 10'd7;
  assign mem[6002] = 10'd8;
  assign mem[6003] = 10'd9;
  assign mem[6004] = 10'd10;
  assign mem[6005] = 10'd11;
  assign mem[6006] = 10'd12;
  assign mem[6007] = 10'd13;
  assign mem[6008] = 10'd14;
  assign mem[6009] = 10'd15;
  assign mem[6010] = 10'd5;
  assign mem[6011] = 10'd6;
  assign mem[6012] = 10'd7;
  assign mem[6013] = 10'd8;
  assign mem[6014] = 10'd9;
  assign mem[6015] = 10'd10;
  assign mem[6016] = 10'd11;
  assign mem[6017] = 10'd12;
  assign mem[6018] = 10'd13;
  assign mem[6019] = 10'd14;
  assign mem[6020] = 10'd4;
  assign mem[6021] = 10'd5;
  assign mem[6022] = 10'd6;
  assign mem[6023] = 10'd7;
  assign mem[6024] = 10'd8;
  assign mem[6025] = 10'd9;
  assign mem[6026] = 10'd10;
  assign mem[6027] = 10'd11;
  assign mem[6028] = 10'd12;
  assign mem[6029] = 10'd13;
  assign mem[6030] = 10'd3;
  assign mem[6031] = 10'd4;
  assign mem[6032] = 10'd5;
  assign mem[6033] = 10'd6;
  assign mem[6034] = 10'd7;
  assign mem[6035] = 10'd8;
  assign mem[6036] = 10'd9;
  assign mem[6037] = 10'd10;
  assign mem[6038] = 10'd11;
  assign mem[6039] = 10'd12;
  assign mem[6040] = 10'd2;
  assign mem[6041] = 10'd3;
  assign mem[6042] = 10'd4;
  assign mem[6043] = 10'd5;
  assign mem[6044] = 10'd6;
  assign mem[6045] = 10'd7;
  assign mem[6046] = 10'd8;
  assign mem[6047] = 10'd9;
  assign mem[6048] = 10'd10;
  assign mem[6049] = 10'd11;
  assign mem[6050] = 10'd1;
  assign mem[6051] = 10'd2;
  assign mem[6052] = 10'd3;
  assign mem[6053] = 10'd4;
  assign mem[6054] = 10'd5;
  assign mem[6055] = 10'd6;
  assign mem[6056] = 10'd7;
  assign mem[6057] = 10'd8;
  assign mem[6058] = 10'd9;
  assign mem[6059] = 10'd10;
  assign mem[6060] = 10'd0;
  assign mem[6061] = 10'd1;
  assign mem[6062] = 10'd2;
  assign mem[6063] = 10'd3;
  assign mem[6064] = 10'd4;
  assign mem[6065] = 10'd5;
  assign mem[6066] = 10'd6;
  assign mem[6067] = 10'd7;
  assign mem[6068] = 10'd8;
  assign mem[6069] = 10'd9;
  assign mem[6070] = 10'd1;
  assign mem[6071] = 10'd2;
  assign mem[6072] = 10'd3;
  assign mem[6073] = 10'd4;
  assign mem[6074] = 10'd5;
  assign mem[6075] = 10'd6;
  assign mem[6076] = 10'd7;
  assign mem[6077] = 10'd8;
  assign mem[6078] = 10'd9;
  assign mem[6079] = 10'd10;
  assign mem[6080] = 10'd2;
  assign mem[6081] = 10'd3;
  assign mem[6082] = 10'd4;
  assign mem[6083] = 10'd5;
  assign mem[6084] = 10'd6;
  assign mem[6085] = 10'd7;
  assign mem[6086] = 10'd8;
  assign mem[6087] = 10'd9;
  assign mem[6088] = 10'd10;
  assign mem[6089] = 10'd11;
  assign mem[6090] = 10'd3;
  assign mem[6091] = 10'd4;
  assign mem[6092] = 10'd5;
  assign mem[6093] = 10'd6;
  assign mem[6094] = 10'd7;
  assign mem[6095] = 10'd8;
  assign mem[6096] = 10'd9;
  assign mem[6097] = 10'd10;
  assign mem[6098] = 10'd11;
  assign mem[6099] = 10'd12;
  assign mem[6100] = 10'd7;
  assign mem[6101] = 10'd6;
  assign mem[6102] = 10'd7;
  assign mem[6103] = 10'd8;
  assign mem[6104] = 10'd9;
  assign mem[6105] = 10'd10;
  assign mem[6106] = 10'd11;
  assign mem[6107] = 10'd12;
  assign mem[6108] = 10'd13;
  assign mem[6109] = 10'd14;
  assign mem[6110] = 10'd6;
  assign mem[6111] = 10'd5;
  assign mem[6112] = 10'd6;
  assign mem[6113] = 10'd7;
  assign mem[6114] = 10'd8;
  assign mem[6115] = 10'd9;
  assign mem[6116] = 10'd10;
  assign mem[6117] = 10'd11;
  assign mem[6118] = 10'd12;
  assign mem[6119] = 10'd13;
  assign mem[6120] = 10'd5;
  assign mem[6121] = 10'd4;
  assign mem[6122] = 10'd5;
  assign mem[6123] = 10'd6;
  assign mem[6124] = 10'd7;
  assign mem[6125] = 10'd8;
  assign mem[6126] = 10'd9;
  assign mem[6127] = 10'd10;
  assign mem[6128] = 10'd11;
  assign mem[6129] = 10'd12;
  assign mem[6130] = 10'd4;
  assign mem[6131] = 10'd3;
  assign mem[6132] = 10'd4;
  assign mem[6133] = 10'd5;
  assign mem[6134] = 10'd6;
  assign mem[6135] = 10'd7;
  assign mem[6136] = 10'd8;
  assign mem[6137] = 10'd9;
  assign mem[6138] = 10'd10;
  assign mem[6139] = 10'd11;
  assign mem[6140] = 10'd3;
  assign mem[6141] = 10'd2;
  assign mem[6142] = 10'd3;
  assign mem[6143] = 10'd4;
  assign mem[6144] = 10'd5;
  assign mem[6145] = 10'd6;
  assign mem[6146] = 10'd7;
  assign mem[6147] = 10'd8;
  assign mem[6148] = 10'd9;
  assign mem[6149] = 10'd10;
  assign mem[6150] = 10'd2;
  assign mem[6151] = 10'd1;
  assign mem[6152] = 10'd2;
  assign mem[6153] = 10'd3;
  assign mem[6154] = 10'd4;
  assign mem[6155] = 10'd5;
  assign mem[6156] = 10'd6;
  assign mem[6157] = 10'd7;
  assign mem[6158] = 10'd8;
  assign mem[6159] = 10'd9;
  assign mem[6160] = 10'd1;
  assign mem[6161] = 10'd0;
  assign mem[6162] = 10'd1;
  assign mem[6163] = 10'd2;
  assign mem[6164] = 10'd3;
  assign mem[6165] = 10'd4;
  assign mem[6166] = 10'd5;
  assign mem[6167] = 10'd6;
  assign mem[6168] = 10'd7;
  assign mem[6169] = 10'd8;
  assign mem[6170] = 10'd2;
  assign mem[6171] = 10'd1;
  assign mem[6172] = 10'd2;
  assign mem[6173] = 10'd3;
  assign mem[6174] = 10'd4;
  assign mem[6175] = 10'd5;
  assign mem[6176] = 10'd6;
  assign mem[6177] = 10'd7;
  assign mem[6178] = 10'd8;
  assign mem[6179] = 10'd9;
  assign mem[6180] = 10'd3;
  assign mem[6181] = 10'd2;
  assign mem[6182] = 10'd3;
  assign mem[6183] = 10'd4;
  assign mem[6184] = 10'd5;
  assign mem[6185] = 10'd6;
  assign mem[6186] = 10'd7;
  assign mem[6187] = 10'd8;
  assign mem[6188] = 10'd9;
  assign mem[6189] = 10'd10;
  assign mem[6190] = 10'd4;
  assign mem[6191] = 10'd3;
  assign mem[6192] = 10'd4;
  assign mem[6193] = 10'd5;
  assign mem[6194] = 10'd6;
  assign mem[6195] = 10'd7;
  assign mem[6196] = 10'd8;
  assign mem[6197] = 10'd9;
  assign mem[6198] = 10'd10;
  assign mem[6199] = 10'd11;
  assign mem[6200] = 10'd8;
  assign mem[6201] = 10'd7;
  assign mem[6202] = 10'd6;
  assign mem[6203] = 10'd7;
  assign mem[6204] = 10'd8;
  assign mem[6205] = 10'd9;
  assign mem[6206] = 10'd10;
  assign mem[6207] = 10'd11;
  assign mem[6208] = 10'd12;
  assign mem[6209] = 10'd13;
  assign mem[6210] = 10'd7;
  assign mem[6211] = 10'd6;
  assign mem[6212] = 10'd5;
  assign mem[6213] = 10'd6;
  assign mem[6214] = 10'd7;
  assign mem[6215] = 10'd8;
  assign mem[6216] = 10'd9;
  assign mem[6217] = 10'd10;
  assign mem[6218] = 10'd11;
  assign mem[6219] = 10'd12;
  assign mem[6220] = 10'd6;
  assign mem[6221] = 10'd5;
  assign mem[6222] = 10'd4;
  assign mem[6223] = 10'd5;
  assign mem[6224] = 10'd6;
  assign mem[6225] = 10'd7;
  assign mem[6226] = 10'd8;
  assign mem[6227] = 10'd9;
  assign mem[6228] = 10'd10;
  assign mem[6229] = 10'd11;
  assign mem[6230] = 10'd5;
  assign mem[6231] = 10'd4;
  assign mem[6232] = 10'd3;
  assign mem[6233] = 10'd4;
  assign mem[6234] = 10'd5;
  assign mem[6235] = 10'd6;
  assign mem[6236] = 10'd7;
  assign mem[6237] = 10'd8;
  assign mem[6238] = 10'd9;
  assign mem[6239] = 10'd10;
  assign mem[6240] = 10'd4;
  assign mem[6241] = 10'd3;
  assign mem[6242] = 10'd2;
  assign mem[6243] = 10'd3;
  assign mem[6244] = 10'd4;
  assign mem[6245] = 10'd5;
  assign mem[6246] = 10'd6;
  assign mem[6247] = 10'd7;
  assign mem[6248] = 10'd8;
  assign mem[6249] = 10'd9;
  assign mem[6250] = 10'd3;
  assign mem[6251] = 10'd2;
  assign mem[6252] = 10'd1;
  assign mem[6253] = 10'd2;
  assign mem[6254] = 10'd3;
  assign mem[6255] = 10'd4;
  assign mem[6256] = 10'd5;
  assign mem[6257] = 10'd6;
  assign mem[6258] = 10'd7;
  assign mem[6259] = 10'd8;
  assign mem[6260] = 10'd2;
  assign mem[6261] = 10'd1;
  assign mem[6262] = 10'd0;
  assign mem[6263] = 10'd1;
  assign mem[6264] = 10'd2;
  assign mem[6265] = 10'd3;
  assign mem[6266] = 10'd4;
  assign mem[6267] = 10'd5;
  assign mem[6268] = 10'd6;
  assign mem[6269] = 10'd7;
  assign mem[6270] = 10'd3;
  assign mem[6271] = 10'd2;
  assign mem[6272] = 10'd1;
  assign mem[6273] = 10'd2;
  assign mem[6274] = 10'd3;
  assign mem[6275] = 10'd4;
  assign mem[6276] = 10'd5;
  assign mem[6277] = 10'd6;
  assign mem[6278] = 10'd7;
  assign mem[6279] = 10'd8;
  assign mem[6280] = 10'd4;
  assign mem[6281] = 10'd3;
  assign mem[6282] = 10'd2;
  assign mem[6283] = 10'd3;
  assign mem[6284] = 10'd4;
  assign mem[6285] = 10'd5;
  assign mem[6286] = 10'd6;
  assign mem[6287] = 10'd7;
  assign mem[6288] = 10'd8;
  assign mem[6289] = 10'd9;
  assign mem[6290] = 10'd5;
  assign mem[6291] = 10'd4;
  assign mem[6292] = 10'd3;
  assign mem[6293] = 10'd4;
  assign mem[6294] = 10'd5;
  assign mem[6295] = 10'd6;
  assign mem[6296] = 10'd7;
  assign mem[6297] = 10'd8;
  assign mem[6298] = 10'd9;
  assign mem[6299] = 10'd10;
  assign mem[6300] = 10'd9;
  assign mem[6301] = 10'd8;
  assign mem[6302] = 10'd7;
  assign mem[6303] = 10'd6;
  assign mem[6304] = 10'd7;
  assign mem[6305] = 10'd8;
  assign mem[6306] = 10'd9;
  assign mem[6307] = 10'd10;
  assign mem[6308] = 10'd11;
  assign mem[6309] = 10'd12;
  assign mem[6310] = 10'd8;
  assign mem[6311] = 10'd7;
  assign mem[6312] = 10'd6;
  assign mem[6313] = 10'd5;
  assign mem[6314] = 10'd6;
  assign mem[6315] = 10'd7;
  assign mem[6316] = 10'd8;
  assign mem[6317] = 10'd9;
  assign mem[6318] = 10'd10;
  assign mem[6319] = 10'd11;
  assign mem[6320] = 10'd7;
  assign mem[6321] = 10'd6;
  assign mem[6322] = 10'd5;
  assign mem[6323] = 10'd4;
  assign mem[6324] = 10'd5;
  assign mem[6325] = 10'd6;
  assign mem[6326] = 10'd7;
  assign mem[6327] = 10'd8;
  assign mem[6328] = 10'd9;
  assign mem[6329] = 10'd10;
  assign mem[6330] = 10'd6;
  assign mem[6331] = 10'd5;
  assign mem[6332] = 10'd4;
  assign mem[6333] = 10'd3;
  assign mem[6334] = 10'd4;
  assign mem[6335] = 10'd5;
  assign mem[6336] = 10'd6;
  assign mem[6337] = 10'd7;
  assign mem[6338] = 10'd8;
  assign mem[6339] = 10'd9;
  assign mem[6340] = 10'd5;
  assign mem[6341] = 10'd4;
  assign mem[6342] = 10'd3;
  assign mem[6343] = 10'd2;
  assign mem[6344] = 10'd3;
  assign mem[6345] = 10'd4;
  assign mem[6346] = 10'd5;
  assign mem[6347] = 10'd6;
  assign mem[6348] = 10'd7;
  assign mem[6349] = 10'd8;
  assign mem[6350] = 10'd4;
  assign mem[6351] = 10'd3;
  assign mem[6352] = 10'd2;
  assign mem[6353] = 10'd1;
  assign mem[6354] = 10'd2;
  assign mem[6355] = 10'd3;
  assign mem[6356] = 10'd4;
  assign mem[6357] = 10'd5;
  assign mem[6358] = 10'd6;
  assign mem[6359] = 10'd7;
  assign mem[6360] = 10'd3;
  assign mem[6361] = 10'd2;
  assign mem[6362] = 10'd1;
  assign mem[6363] = 10'd0;
  assign mem[6364] = 10'd1;
  assign mem[6365] = 10'd2;
  assign mem[6366] = 10'd3;
  assign mem[6367] = 10'd4;
  assign mem[6368] = 10'd5;
  assign mem[6369] = 10'd6;
  assign mem[6370] = 10'd4;
  assign mem[6371] = 10'd3;
  assign mem[6372] = 10'd2;
  assign mem[6373] = 10'd1;
  assign mem[6374] = 10'd2;
  assign mem[6375] = 10'd3;
  assign mem[6376] = 10'd4;
  assign mem[6377] = 10'd5;
  assign mem[6378] = 10'd6;
  assign mem[6379] = 10'd7;
  assign mem[6380] = 10'd5;
  assign mem[6381] = 10'd4;
  assign mem[6382] = 10'd3;
  assign mem[6383] = 10'd2;
  assign mem[6384] = 10'd3;
  assign mem[6385] = 10'd4;
  assign mem[6386] = 10'd5;
  assign mem[6387] = 10'd6;
  assign mem[6388] = 10'd7;
  assign mem[6389] = 10'd8;
  assign mem[6390] = 10'd6;
  assign mem[6391] = 10'd5;
  assign mem[6392] = 10'd4;
  assign mem[6393] = 10'd3;
  assign mem[6394] = 10'd4;
  assign mem[6395] = 10'd5;
  assign mem[6396] = 10'd6;
  assign mem[6397] = 10'd7;
  assign mem[6398] = 10'd8;
  assign mem[6399] = 10'd9;
  assign mem[6400] = 10'd10;
  assign mem[6401] = 10'd9;
  assign mem[6402] = 10'd8;
  assign mem[6403] = 10'd7;
  assign mem[6404] = 10'd6;
  assign mem[6405] = 10'd7;
  assign mem[6406] = 10'd8;
  assign mem[6407] = 10'd9;
  assign mem[6408] = 10'd10;
  assign mem[6409] = 10'd11;
  assign mem[6410] = 10'd9;
  assign mem[6411] = 10'd8;
  assign mem[6412] = 10'd7;
  assign mem[6413] = 10'd6;
  assign mem[6414] = 10'd5;
  assign mem[6415] = 10'd6;
  assign mem[6416] = 10'd7;
  assign mem[6417] = 10'd8;
  assign mem[6418] = 10'd9;
  assign mem[6419] = 10'd10;
  assign mem[6420] = 10'd8;
  assign mem[6421] = 10'd7;
  assign mem[6422] = 10'd6;
  assign mem[6423] = 10'd5;
  assign mem[6424] = 10'd4;
  assign mem[6425] = 10'd5;
  assign mem[6426] = 10'd6;
  assign mem[6427] = 10'd7;
  assign mem[6428] = 10'd8;
  assign mem[6429] = 10'd9;
  assign mem[6430] = 10'd7;
  assign mem[6431] = 10'd6;
  assign mem[6432] = 10'd5;
  assign mem[6433] = 10'd4;
  assign mem[6434] = 10'd3;
  assign mem[6435] = 10'd4;
  assign mem[6436] = 10'd5;
  assign mem[6437] = 10'd6;
  assign mem[6438] = 10'd7;
  assign mem[6439] = 10'd8;
  assign mem[6440] = 10'd6;
  assign mem[6441] = 10'd5;
  assign mem[6442] = 10'd4;
  assign mem[6443] = 10'd3;
  assign mem[6444] = 10'd2;
  assign mem[6445] = 10'd3;
  assign mem[6446] = 10'd4;
  assign mem[6447] = 10'd5;
  assign mem[6448] = 10'd6;
  assign mem[6449] = 10'd7;
  assign mem[6450] = 10'd5;
  assign mem[6451] = 10'd4;
  assign mem[6452] = 10'd3;
  assign mem[6453] = 10'd2;
  assign mem[6454] = 10'd1;
  assign mem[6455] = 10'd2;
  assign mem[6456] = 10'd3;
  assign mem[6457] = 10'd4;
  assign mem[6458] = 10'd5;
  assign mem[6459] = 10'd6;
  assign mem[6460] = 10'd4;
  assign mem[6461] = 10'd3;
  assign mem[6462] = 10'd2;
  assign mem[6463] = 10'd1;
  assign mem[6464] = 10'd0;
  assign mem[6465] = 10'd1;
  assign mem[6466] = 10'd2;
  assign mem[6467] = 10'd3;
  assign mem[6468] = 10'd4;
  assign mem[6469] = 10'd5;
  assign mem[6470] = 10'd5;
  assign mem[6471] = 10'd4;
  assign mem[6472] = 10'd3;
  assign mem[6473] = 10'd2;
  assign mem[6474] = 10'd1;
  assign mem[6475] = 10'd2;
  assign mem[6476] = 10'd3;
  assign mem[6477] = 10'd4;
  assign mem[6478] = 10'd5;
  assign mem[6479] = 10'd6;
  assign mem[6480] = 10'd6;
  assign mem[6481] = 10'd5;
  assign mem[6482] = 10'd4;
  assign mem[6483] = 10'd3;
  assign mem[6484] = 10'd2;
  assign mem[6485] = 10'd3;
  assign mem[6486] = 10'd4;
  assign mem[6487] = 10'd5;
  assign mem[6488] = 10'd6;
  assign mem[6489] = 10'd7;
  assign mem[6490] = 10'd7;
  assign mem[6491] = 10'd6;
  assign mem[6492] = 10'd5;
  assign mem[6493] = 10'd4;
  assign mem[6494] = 10'd3;
  assign mem[6495] = 10'd4;
  assign mem[6496] = 10'd5;
  assign mem[6497] = 10'd6;
  assign mem[6498] = 10'd7;
  assign mem[6499] = 10'd8;
  assign mem[6500] = 10'd11;
  assign mem[6501] = 10'd10;
  assign mem[6502] = 10'd9;
  assign mem[6503] = 10'd8;
  assign mem[6504] = 10'd7;
  assign mem[6505] = 10'd6;
  assign mem[6506] = 10'd7;
  assign mem[6507] = 10'd8;
  assign mem[6508] = 10'd9;
  assign mem[6509] = 10'd10;
  assign mem[6510] = 10'd10;
  assign mem[6511] = 10'd9;
  assign mem[6512] = 10'd8;
  assign mem[6513] = 10'd7;
  assign mem[6514] = 10'd6;
  assign mem[6515] = 10'd5;
  assign mem[6516] = 10'd6;
  assign mem[6517] = 10'd7;
  assign mem[6518] = 10'd8;
  assign mem[6519] = 10'd9;
  assign mem[6520] = 10'd9;
  assign mem[6521] = 10'd8;
  assign mem[6522] = 10'd7;
  assign mem[6523] = 10'd6;
  assign mem[6524] = 10'd5;
  assign mem[6525] = 10'd4;
  assign mem[6526] = 10'd5;
  assign mem[6527] = 10'd6;
  assign mem[6528] = 10'd7;
  assign mem[6529] = 10'd8;
  assign mem[6530] = 10'd8;
  assign mem[6531] = 10'd7;
  assign mem[6532] = 10'd6;
  assign mem[6533] = 10'd5;
  assign mem[6534] = 10'd4;
  assign mem[6535] = 10'd3;
  assign mem[6536] = 10'd4;
  assign mem[6537] = 10'd5;
  assign mem[6538] = 10'd6;
  assign mem[6539] = 10'd7;
  assign mem[6540] = 10'd7;
  assign mem[6541] = 10'd6;
  assign mem[6542] = 10'd5;
  assign mem[6543] = 10'd4;
  assign mem[6544] = 10'd3;
  assign mem[6545] = 10'd2;
  assign mem[6546] = 10'd3;
  assign mem[6547] = 10'd4;
  assign mem[6548] = 10'd5;
  assign mem[6549] = 10'd6;
  assign mem[6550] = 10'd6;
  assign mem[6551] = 10'd5;
  assign mem[6552] = 10'd4;
  assign mem[6553] = 10'd3;
  assign mem[6554] = 10'd2;
  assign mem[6555] = 10'd1;
  assign mem[6556] = 10'd2;
  assign mem[6557] = 10'd3;
  assign mem[6558] = 10'd4;
  assign mem[6559] = 10'd5;
  assign mem[6560] = 10'd5;
  assign mem[6561] = 10'd4;
  assign mem[6562] = 10'd3;
  assign mem[6563] = 10'd2;
  assign mem[6564] = 10'd1;
  assign mem[6565] = 10'd0;
  assign mem[6566] = 10'd1;
  assign mem[6567] = 10'd2;
  assign mem[6568] = 10'd3;
  assign mem[6569] = 10'd4;
  assign mem[6570] = 10'd6;
  assign mem[6571] = 10'd5;
  assign mem[6572] = 10'd4;
  assign mem[6573] = 10'd3;
  assign mem[6574] = 10'd2;
  assign mem[6575] = 10'd1;
  assign mem[6576] = 10'd2;
  assign mem[6577] = 10'd3;
  assign mem[6578] = 10'd4;
  assign mem[6579] = 10'd5;
  assign mem[6580] = 10'd7;
  assign mem[6581] = 10'd6;
  assign mem[6582] = 10'd5;
  assign mem[6583] = 10'd4;
  assign mem[6584] = 10'd3;
  assign mem[6585] = 10'd2;
  assign mem[6586] = 10'd3;
  assign mem[6587] = 10'd4;
  assign mem[6588] = 10'd5;
  assign mem[6589] = 10'd6;
  assign mem[6590] = 10'd8;
  assign mem[6591] = 10'd7;
  assign mem[6592] = 10'd6;
  assign mem[6593] = 10'd5;
  assign mem[6594] = 10'd4;
  assign mem[6595] = 10'd3;
  assign mem[6596] = 10'd4;
  assign mem[6597] = 10'd5;
  assign mem[6598] = 10'd6;
  assign mem[6599] = 10'd7;
  assign mem[6600] = 10'd12;
  assign mem[6601] = 10'd11;
  assign mem[6602] = 10'd10;
  assign mem[6603] = 10'd9;
  assign mem[6604] = 10'd8;
  assign mem[6605] = 10'd7;
  assign mem[6606] = 10'd6;
  assign mem[6607] = 10'd7;
  assign mem[6608] = 10'd8;
  assign mem[6609] = 10'd9;
  assign mem[6610] = 10'd11;
  assign mem[6611] = 10'd10;
  assign mem[6612] = 10'd9;
  assign mem[6613] = 10'd8;
  assign mem[6614] = 10'd7;
  assign mem[6615] = 10'd6;
  assign mem[6616] = 10'd5;
  assign mem[6617] = 10'd6;
  assign mem[6618] = 10'd7;
  assign mem[6619] = 10'd8;
  assign mem[6620] = 10'd10;
  assign mem[6621] = 10'd9;
  assign mem[6622] = 10'd8;
  assign mem[6623] = 10'd7;
  assign mem[6624] = 10'd6;
  assign mem[6625] = 10'd5;
  assign mem[6626] = 10'd4;
  assign mem[6627] = 10'd5;
  assign mem[6628] = 10'd6;
  assign mem[6629] = 10'd7;
  assign mem[6630] = 10'd9;
  assign mem[6631] = 10'd8;
  assign mem[6632] = 10'd7;
  assign mem[6633] = 10'd6;
  assign mem[6634] = 10'd5;
  assign mem[6635] = 10'd4;
  assign mem[6636] = 10'd3;
  assign mem[6637] = 10'd4;
  assign mem[6638] = 10'd5;
  assign mem[6639] = 10'd6;
  assign mem[6640] = 10'd8;
  assign mem[6641] = 10'd7;
  assign mem[6642] = 10'd6;
  assign mem[6643] = 10'd5;
  assign mem[6644] = 10'd4;
  assign mem[6645] = 10'd3;
  assign mem[6646] = 10'd2;
  assign mem[6647] = 10'd3;
  assign mem[6648] = 10'd4;
  assign mem[6649] = 10'd5;
  assign mem[6650] = 10'd7;
  assign mem[6651] = 10'd6;
  assign mem[6652] = 10'd5;
  assign mem[6653] = 10'd4;
  assign mem[6654] = 10'd3;
  assign mem[6655] = 10'd2;
  assign mem[6656] = 10'd1;
  assign mem[6657] = 10'd2;
  assign mem[6658] = 10'd3;
  assign mem[6659] = 10'd4;
  assign mem[6660] = 10'd6;
  assign mem[6661] = 10'd5;
  assign mem[6662] = 10'd4;
  assign mem[6663] = 10'd3;
  assign mem[6664] = 10'd2;
  assign mem[6665] = 10'd1;
  assign mem[6666] = 10'd0;
  assign mem[6667] = 10'd1;
  assign mem[6668] = 10'd2;
  assign mem[6669] = 10'd3;
  assign mem[6670] = 10'd7;
  assign mem[6671] = 10'd6;
  assign mem[6672] = 10'd5;
  assign mem[6673] = 10'd4;
  assign mem[6674] = 10'd3;
  assign mem[6675] = 10'd2;
  assign mem[6676] = 10'd1;
  assign mem[6677] = 10'd2;
  assign mem[6678] = 10'd3;
  assign mem[6679] = 10'd4;
  assign mem[6680] = 10'd8;
  assign mem[6681] = 10'd7;
  assign mem[6682] = 10'd6;
  assign mem[6683] = 10'd5;
  assign mem[6684] = 10'd4;
  assign mem[6685] = 10'd3;
  assign mem[6686] = 10'd2;
  assign mem[6687] = 10'd3;
  assign mem[6688] = 10'd4;
  assign mem[6689] = 10'd5;
  assign mem[6690] = 10'd9;
  assign mem[6691] = 10'd8;
  assign mem[6692] = 10'd7;
  assign mem[6693] = 10'd6;
  assign mem[6694] = 10'd5;
  assign mem[6695] = 10'd4;
  assign mem[6696] = 10'd3;
  assign mem[6697] = 10'd4;
  assign mem[6698] = 10'd5;
  assign mem[6699] = 10'd6;
  assign mem[6700] = 10'd13;
  assign mem[6701] = 10'd12;
  assign mem[6702] = 10'd11;
  assign mem[6703] = 10'd10;
  assign mem[6704] = 10'd9;
  assign mem[6705] = 10'd8;
  assign mem[6706] = 10'd7;
  assign mem[6707] = 10'd6;
  assign mem[6708] = 10'd7;
  assign mem[6709] = 10'd8;
  assign mem[6710] = 10'd12;
  assign mem[6711] = 10'd11;
  assign mem[6712] = 10'd10;
  assign mem[6713] = 10'd9;
  assign mem[6714] = 10'd8;
  assign mem[6715] = 10'd7;
  assign mem[6716] = 10'd6;
  assign mem[6717] = 10'd5;
  assign mem[6718] = 10'd6;
  assign mem[6719] = 10'd7;
  assign mem[6720] = 10'd11;
  assign mem[6721] = 10'd10;
  assign mem[6722] = 10'd9;
  assign mem[6723] = 10'd8;
  assign mem[6724] = 10'd7;
  assign mem[6725] = 10'd6;
  assign mem[6726] = 10'd5;
  assign mem[6727] = 10'd4;
  assign mem[6728] = 10'd5;
  assign mem[6729] = 10'd6;
  assign mem[6730] = 10'd10;
  assign mem[6731] = 10'd9;
  assign mem[6732] = 10'd8;
  assign mem[6733] = 10'd7;
  assign mem[6734] = 10'd6;
  assign mem[6735] = 10'd5;
  assign mem[6736] = 10'd4;
  assign mem[6737] = 10'd3;
  assign mem[6738] = 10'd4;
  assign mem[6739] = 10'd5;
  assign mem[6740] = 10'd9;
  assign mem[6741] = 10'd8;
  assign mem[6742] = 10'd7;
  assign mem[6743] = 10'd6;
  assign mem[6744] = 10'd5;
  assign mem[6745] = 10'd4;
  assign mem[6746] = 10'd3;
  assign mem[6747] = 10'd2;
  assign mem[6748] = 10'd3;
  assign mem[6749] = 10'd4;
  assign mem[6750] = 10'd8;
  assign mem[6751] = 10'd7;
  assign mem[6752] = 10'd6;
  assign mem[6753] = 10'd5;
  assign mem[6754] = 10'd4;
  assign mem[6755] = 10'd3;
  assign mem[6756] = 10'd2;
  assign mem[6757] = 10'd1;
  assign mem[6758] = 10'd2;
  assign mem[6759] = 10'd3;
  assign mem[6760] = 10'd7;
  assign mem[6761] = 10'd6;
  assign mem[6762] = 10'd5;
  assign mem[6763] = 10'd4;
  assign mem[6764] = 10'd3;
  assign mem[6765] = 10'd2;
  assign mem[6766] = 10'd1;
  assign mem[6767] = 10'd0;
  assign mem[6768] = 10'd1;
  assign mem[6769] = 10'd2;
  assign mem[6770] = 10'd8;
  assign mem[6771] = 10'd7;
  assign mem[6772] = 10'd6;
  assign mem[6773] = 10'd5;
  assign mem[6774] = 10'd4;
  assign mem[6775] = 10'd3;
  assign mem[6776] = 10'd2;
  assign mem[6777] = 10'd1;
  assign mem[6778] = 10'd2;
  assign mem[6779] = 10'd3;
  assign mem[6780] = 10'd9;
  assign mem[6781] = 10'd8;
  assign mem[6782] = 10'd7;
  assign mem[6783] = 10'd6;
  assign mem[6784] = 10'd5;
  assign mem[6785] = 10'd4;
  assign mem[6786] = 10'd3;
  assign mem[6787] = 10'd2;
  assign mem[6788] = 10'd3;
  assign mem[6789] = 10'd4;
  assign mem[6790] = 10'd10;
  assign mem[6791] = 10'd9;
  assign mem[6792] = 10'd8;
  assign mem[6793] = 10'd7;
  assign mem[6794] = 10'd6;
  assign mem[6795] = 10'd5;
  assign mem[6796] = 10'd4;
  assign mem[6797] = 10'd3;
  assign mem[6798] = 10'd4;
  assign mem[6799] = 10'd5;
  assign mem[6800] = 10'd14;
  assign mem[6801] = 10'd13;
  assign mem[6802] = 10'd12;
  assign mem[6803] = 10'd11;
  assign mem[6804] = 10'd10;
  assign mem[6805] = 10'd9;
  assign mem[6806] = 10'd8;
  assign mem[6807] = 10'd7;
  assign mem[6808] = 10'd6;
  assign mem[6809] = 10'd7;
  assign mem[6810] = 10'd13;
  assign mem[6811] = 10'd12;
  assign mem[6812] = 10'd11;
  assign mem[6813] = 10'd10;
  assign mem[6814] = 10'd9;
  assign mem[6815] = 10'd8;
  assign mem[6816] = 10'd7;
  assign mem[6817] = 10'd6;
  assign mem[6818] = 10'd5;
  assign mem[6819] = 10'd6;
  assign mem[6820] = 10'd12;
  assign mem[6821] = 10'd11;
  assign mem[6822] = 10'd10;
  assign mem[6823] = 10'd9;
  assign mem[6824] = 10'd8;
  assign mem[6825] = 10'd7;
  assign mem[6826] = 10'd6;
  assign mem[6827] = 10'd5;
  assign mem[6828] = 10'd4;
  assign mem[6829] = 10'd5;
  assign mem[6830] = 10'd11;
  assign mem[6831] = 10'd10;
  assign mem[6832] = 10'd9;
  assign mem[6833] = 10'd8;
  assign mem[6834] = 10'd7;
  assign mem[6835] = 10'd6;
  assign mem[6836] = 10'd5;
  assign mem[6837] = 10'd4;
  assign mem[6838] = 10'd3;
  assign mem[6839] = 10'd4;
  assign mem[6840] = 10'd10;
  assign mem[6841] = 10'd9;
  assign mem[6842] = 10'd8;
  assign mem[6843] = 10'd7;
  assign mem[6844] = 10'd6;
  assign mem[6845] = 10'd5;
  assign mem[6846] = 10'd4;
  assign mem[6847] = 10'd3;
  assign mem[6848] = 10'd2;
  assign mem[6849] = 10'd3;
  assign mem[6850] = 10'd9;
  assign mem[6851] = 10'd8;
  assign mem[6852] = 10'd7;
  assign mem[6853] = 10'd6;
  assign mem[6854] = 10'd5;
  assign mem[6855] = 10'd4;
  assign mem[6856] = 10'd3;
  assign mem[6857] = 10'd2;
  assign mem[6858] = 10'd1;
  assign mem[6859] = 10'd2;
  assign mem[6860] = 10'd8;
  assign mem[6861] = 10'd7;
  assign mem[6862] = 10'd6;
  assign mem[6863] = 10'd5;
  assign mem[6864] = 10'd4;
  assign mem[6865] = 10'd3;
  assign mem[6866] = 10'd2;
  assign mem[6867] = 10'd1;
  assign mem[6868] = 10'd0;
  assign mem[6869] = 10'd1;
  assign mem[6870] = 10'd9;
  assign mem[6871] = 10'd8;
  assign mem[6872] = 10'd7;
  assign mem[6873] = 10'd6;
  assign mem[6874] = 10'd5;
  assign mem[6875] = 10'd4;
  assign mem[6876] = 10'd3;
  assign mem[6877] = 10'd2;
  assign mem[6878] = 10'd1;
  assign mem[6879] = 10'd2;
  assign mem[6880] = 10'd10;
  assign mem[6881] = 10'd9;
  assign mem[6882] = 10'd8;
  assign mem[6883] = 10'd7;
  assign mem[6884] = 10'd6;
  assign mem[6885] = 10'd5;
  assign mem[6886] = 10'd4;
  assign mem[6887] = 10'd3;
  assign mem[6888] = 10'd2;
  assign mem[6889] = 10'd3;
  assign mem[6890] = 10'd11;
  assign mem[6891] = 10'd10;
  assign mem[6892] = 10'd9;
  assign mem[6893] = 10'd8;
  assign mem[6894] = 10'd7;
  assign mem[6895] = 10'd6;
  assign mem[6896] = 10'd5;
  assign mem[6897] = 10'd4;
  assign mem[6898] = 10'd3;
  assign mem[6899] = 10'd4;
  assign mem[6900] = 10'd15;
  assign mem[6901] = 10'd14;
  assign mem[6902] = 10'd13;
  assign mem[6903] = 10'd12;
  assign mem[6904] = 10'd11;
  assign mem[6905] = 10'd10;
  assign mem[6906] = 10'd9;
  assign mem[6907] = 10'd8;
  assign mem[6908] = 10'd7;
  assign mem[6909] = 10'd6;
  assign mem[6910] = 10'd14;
  assign mem[6911] = 10'd13;
  assign mem[6912] = 10'd12;
  assign mem[6913] = 10'd11;
  assign mem[6914] = 10'd10;
  assign mem[6915] = 10'd9;
  assign mem[6916] = 10'd8;
  assign mem[6917] = 10'd7;
  assign mem[6918] = 10'd6;
  assign mem[6919] = 10'd5;
  assign mem[6920] = 10'd13;
  assign mem[6921] = 10'd12;
  assign mem[6922] = 10'd11;
  assign mem[6923] = 10'd10;
  assign mem[6924] = 10'd9;
  assign mem[6925] = 10'd8;
  assign mem[6926] = 10'd7;
  assign mem[6927] = 10'd6;
  assign mem[6928] = 10'd5;
  assign mem[6929] = 10'd4;
  assign mem[6930] = 10'd12;
  assign mem[6931] = 10'd11;
  assign mem[6932] = 10'd10;
  assign mem[6933] = 10'd9;
  assign mem[6934] = 10'd8;
  assign mem[6935] = 10'd7;
  assign mem[6936] = 10'd6;
  assign mem[6937] = 10'd5;
  assign mem[6938] = 10'd4;
  assign mem[6939] = 10'd3;
  assign mem[6940] = 10'd11;
  assign mem[6941] = 10'd10;
  assign mem[6942] = 10'd9;
  assign mem[6943] = 10'd8;
  assign mem[6944] = 10'd7;
  assign mem[6945] = 10'd6;
  assign mem[6946] = 10'd5;
  assign mem[6947] = 10'd4;
  assign mem[6948] = 10'd3;
  assign mem[6949] = 10'd2;
  assign mem[6950] = 10'd10;
  assign mem[6951] = 10'd9;
  assign mem[6952] = 10'd8;
  assign mem[6953] = 10'd7;
  assign mem[6954] = 10'd6;
  assign mem[6955] = 10'd5;
  assign mem[6956] = 10'd4;
  assign mem[6957] = 10'd3;
  assign mem[6958] = 10'd2;
  assign mem[6959] = 10'd1;
  assign mem[6960] = 10'd9;
  assign mem[6961] = 10'd8;
  assign mem[6962] = 10'd7;
  assign mem[6963] = 10'd6;
  assign mem[6964] = 10'd5;
  assign mem[6965] = 10'd4;
  assign mem[6966] = 10'd3;
  assign mem[6967] = 10'd2;
  assign mem[6968] = 10'd1;
  assign mem[6969] = 10'd0;
  assign mem[6970] = 10'd10;
  assign mem[6971] = 10'd9;
  assign mem[6972] = 10'd8;
  assign mem[6973] = 10'd7;
  assign mem[6974] = 10'd6;
  assign mem[6975] = 10'd5;
  assign mem[6976] = 10'd4;
  assign mem[6977] = 10'd3;
  assign mem[6978] = 10'd2;
  assign mem[6979] = 10'd1;
  assign mem[6980] = 10'd11;
  assign mem[6981] = 10'd10;
  assign mem[6982] = 10'd9;
  assign mem[6983] = 10'd8;
  assign mem[6984] = 10'd7;
  assign mem[6985] = 10'd6;
  assign mem[6986] = 10'd5;
  assign mem[6987] = 10'd4;
  assign mem[6988] = 10'd3;
  assign mem[6989] = 10'd2;
  assign mem[6990] = 10'd12;
  assign mem[6991] = 10'd11;
  assign mem[6992] = 10'd10;
  assign mem[6993] = 10'd9;
  assign mem[6994] = 10'd8;
  assign mem[6995] = 10'd7;
  assign mem[6996] = 10'd6;
  assign mem[6997] = 10'd5;
  assign mem[6998] = 10'd4;
  assign mem[6999] = 10'd3;
  assign mem[7000] = 10'd7;
  assign mem[7001] = 10'd8;
  assign mem[7002] = 10'd9;
  assign mem[7003] = 10'd10;
  assign mem[7004] = 10'd11;
  assign mem[7005] = 10'd12;
  assign mem[7006] = 10'd13;
  assign mem[7007] = 10'd14;
  assign mem[7008] = 10'd15;
  assign mem[7009] = 10'd16;
  assign mem[7010] = 10'd6;
  assign mem[7011] = 10'd7;
  assign mem[7012] = 10'd8;
  assign mem[7013] = 10'd9;
  assign mem[7014] = 10'd10;
  assign mem[7015] = 10'd11;
  assign mem[7016] = 10'd12;
  assign mem[7017] = 10'd13;
  assign mem[7018] = 10'd14;
  assign mem[7019] = 10'd15;
  assign mem[7020] = 10'd5;
  assign mem[7021] = 10'd6;
  assign mem[7022] = 10'd7;
  assign mem[7023] = 10'd8;
  assign mem[7024] = 10'd9;
  assign mem[7025] = 10'd10;
  assign mem[7026] = 10'd11;
  assign mem[7027] = 10'd12;
  assign mem[7028] = 10'd13;
  assign mem[7029] = 10'd14;
  assign mem[7030] = 10'd4;
  assign mem[7031] = 10'd5;
  assign mem[7032] = 10'd6;
  assign mem[7033] = 10'd7;
  assign mem[7034] = 10'd8;
  assign mem[7035] = 10'd9;
  assign mem[7036] = 10'd10;
  assign mem[7037] = 10'd11;
  assign mem[7038] = 10'd12;
  assign mem[7039] = 10'd13;
  assign mem[7040] = 10'd3;
  assign mem[7041] = 10'd4;
  assign mem[7042] = 10'd5;
  assign mem[7043] = 10'd6;
  assign mem[7044] = 10'd7;
  assign mem[7045] = 10'd8;
  assign mem[7046] = 10'd9;
  assign mem[7047] = 10'd10;
  assign mem[7048] = 10'd11;
  assign mem[7049] = 10'd12;
  assign mem[7050] = 10'd2;
  assign mem[7051] = 10'd3;
  assign mem[7052] = 10'd4;
  assign mem[7053] = 10'd5;
  assign mem[7054] = 10'd6;
  assign mem[7055] = 10'd7;
  assign mem[7056] = 10'd8;
  assign mem[7057] = 10'd9;
  assign mem[7058] = 10'd10;
  assign mem[7059] = 10'd11;
  assign mem[7060] = 10'd1;
  assign mem[7061] = 10'd2;
  assign mem[7062] = 10'd3;
  assign mem[7063] = 10'd4;
  assign mem[7064] = 10'd5;
  assign mem[7065] = 10'd6;
  assign mem[7066] = 10'd7;
  assign mem[7067] = 10'd8;
  assign mem[7068] = 10'd9;
  assign mem[7069] = 10'd10;
  assign mem[7070] = 10'd0;
  assign mem[7071] = 10'd1;
  assign mem[7072] = 10'd2;
  assign mem[7073] = 10'd3;
  assign mem[7074] = 10'd4;
  assign mem[7075] = 10'd5;
  assign mem[7076] = 10'd6;
  assign mem[7077] = 10'd7;
  assign mem[7078] = 10'd8;
  assign mem[7079] = 10'd9;
  assign mem[7080] = 10'd1;
  assign mem[7081] = 10'd2;
  assign mem[7082] = 10'd3;
  assign mem[7083] = 10'd4;
  assign mem[7084] = 10'd5;
  assign mem[7085] = 10'd6;
  assign mem[7086] = 10'd7;
  assign mem[7087] = 10'd8;
  assign mem[7088] = 10'd9;
  assign mem[7089] = 10'd10;
  assign mem[7090] = 10'd2;
  assign mem[7091] = 10'd3;
  assign mem[7092] = 10'd4;
  assign mem[7093] = 10'd5;
  assign mem[7094] = 10'd6;
  assign mem[7095] = 10'd7;
  assign mem[7096] = 10'd8;
  assign mem[7097] = 10'd9;
  assign mem[7098] = 10'd10;
  assign mem[7099] = 10'd11;
  assign mem[7100] = 10'd8;
  assign mem[7101] = 10'd7;
  assign mem[7102] = 10'd8;
  assign mem[7103] = 10'd9;
  assign mem[7104] = 10'd10;
  assign mem[7105] = 10'd11;
  assign mem[7106] = 10'd12;
  assign mem[7107] = 10'd13;
  assign mem[7108] = 10'd14;
  assign mem[7109] = 10'd15;
  assign mem[7110] = 10'd7;
  assign mem[7111] = 10'd6;
  assign mem[7112] = 10'd7;
  assign mem[7113] = 10'd8;
  assign mem[7114] = 10'd9;
  assign mem[7115] = 10'd10;
  assign mem[7116] = 10'd11;
  assign mem[7117] = 10'd12;
  assign mem[7118] = 10'd13;
  assign mem[7119] = 10'd14;
  assign mem[7120] = 10'd6;
  assign mem[7121] = 10'd5;
  assign mem[7122] = 10'd6;
  assign mem[7123] = 10'd7;
  assign mem[7124] = 10'd8;
  assign mem[7125] = 10'd9;
  assign mem[7126] = 10'd10;
  assign mem[7127] = 10'd11;
  assign mem[7128] = 10'd12;
  assign mem[7129] = 10'd13;
  assign mem[7130] = 10'd5;
  assign mem[7131] = 10'd4;
  assign mem[7132] = 10'd5;
  assign mem[7133] = 10'd6;
  assign mem[7134] = 10'd7;
  assign mem[7135] = 10'd8;
  assign mem[7136] = 10'd9;
  assign mem[7137] = 10'd10;
  assign mem[7138] = 10'd11;
  assign mem[7139] = 10'd12;
  assign mem[7140] = 10'd4;
  assign mem[7141] = 10'd3;
  assign mem[7142] = 10'd4;
  assign mem[7143] = 10'd5;
  assign mem[7144] = 10'd6;
  assign mem[7145] = 10'd7;
  assign mem[7146] = 10'd8;
  assign mem[7147] = 10'd9;
  assign mem[7148] = 10'd10;
  assign mem[7149] = 10'd11;
  assign mem[7150] = 10'd3;
  assign mem[7151] = 10'd2;
  assign mem[7152] = 10'd3;
  assign mem[7153] = 10'd4;
  assign mem[7154] = 10'd5;
  assign mem[7155] = 10'd6;
  assign mem[7156] = 10'd7;
  assign mem[7157] = 10'd8;
  assign mem[7158] = 10'd9;
  assign mem[7159] = 10'd10;
  assign mem[7160] = 10'd2;
  assign mem[7161] = 10'd1;
  assign mem[7162] = 10'd2;
  assign mem[7163] = 10'd3;
  assign mem[7164] = 10'd4;
  assign mem[7165] = 10'd5;
  assign mem[7166] = 10'd6;
  assign mem[7167] = 10'd7;
  assign mem[7168] = 10'd8;
  assign mem[7169] = 10'd9;
  assign mem[7170] = 10'd1;
  assign mem[7171] = 10'd0;
  assign mem[7172] = 10'd1;
  assign mem[7173] = 10'd2;
  assign mem[7174] = 10'd3;
  assign mem[7175] = 10'd4;
  assign mem[7176] = 10'd5;
  assign mem[7177] = 10'd6;
  assign mem[7178] = 10'd7;
  assign mem[7179] = 10'd8;
  assign mem[7180] = 10'd2;
  assign mem[7181] = 10'd1;
  assign mem[7182] = 10'd2;
  assign mem[7183] = 10'd3;
  assign mem[7184] = 10'd4;
  assign mem[7185] = 10'd5;
  assign mem[7186] = 10'd6;
  assign mem[7187] = 10'd7;
  assign mem[7188] = 10'd8;
  assign mem[7189] = 10'd9;
  assign mem[7190] = 10'd3;
  assign mem[7191] = 10'd2;
  assign mem[7192] = 10'd3;
  assign mem[7193] = 10'd4;
  assign mem[7194] = 10'd5;
  assign mem[7195] = 10'd6;
  assign mem[7196] = 10'd7;
  assign mem[7197] = 10'd8;
  assign mem[7198] = 10'd9;
  assign mem[7199] = 10'd10;
  assign mem[7200] = 10'd9;
  assign mem[7201] = 10'd8;
  assign mem[7202] = 10'd7;
  assign mem[7203] = 10'd8;
  assign mem[7204] = 10'd9;
  assign mem[7205] = 10'd10;
  assign mem[7206] = 10'd11;
  assign mem[7207] = 10'd12;
  assign mem[7208] = 10'd13;
  assign mem[7209] = 10'd14;
  assign mem[7210] = 10'd8;
  assign mem[7211] = 10'd7;
  assign mem[7212] = 10'd6;
  assign mem[7213] = 10'd7;
  assign mem[7214] = 10'd8;
  assign mem[7215] = 10'd9;
  assign mem[7216] = 10'd10;
  assign mem[7217] = 10'd11;
  assign mem[7218] = 10'd12;
  assign mem[7219] = 10'd13;
  assign mem[7220] = 10'd7;
  assign mem[7221] = 10'd6;
  assign mem[7222] = 10'd5;
  assign mem[7223] = 10'd6;
  assign mem[7224] = 10'd7;
  assign mem[7225] = 10'd8;
  assign mem[7226] = 10'd9;
  assign mem[7227] = 10'd10;
  assign mem[7228] = 10'd11;
  assign mem[7229] = 10'd12;
  assign mem[7230] = 10'd6;
  assign mem[7231] = 10'd5;
  assign mem[7232] = 10'd4;
  assign mem[7233] = 10'd5;
  assign mem[7234] = 10'd6;
  assign mem[7235] = 10'd7;
  assign mem[7236] = 10'd8;
  assign mem[7237] = 10'd9;
  assign mem[7238] = 10'd10;
  assign mem[7239] = 10'd11;
  assign mem[7240] = 10'd5;
  assign mem[7241] = 10'd4;
  assign mem[7242] = 10'd3;
  assign mem[7243] = 10'd4;
  assign mem[7244] = 10'd5;
  assign mem[7245] = 10'd6;
  assign mem[7246] = 10'd7;
  assign mem[7247] = 10'd8;
  assign mem[7248] = 10'd9;
  assign mem[7249] = 10'd10;
  assign mem[7250] = 10'd4;
  assign mem[7251] = 10'd3;
  assign mem[7252] = 10'd2;
  assign mem[7253] = 10'd3;
  assign mem[7254] = 10'd4;
  assign mem[7255] = 10'd5;
  assign mem[7256] = 10'd6;
  assign mem[7257] = 10'd7;
  assign mem[7258] = 10'd8;
  assign mem[7259] = 10'd9;
  assign mem[7260] = 10'd3;
  assign mem[7261] = 10'd2;
  assign mem[7262] = 10'd1;
  assign mem[7263] = 10'd2;
  assign mem[7264] = 10'd3;
  assign mem[7265] = 10'd4;
  assign mem[7266] = 10'd5;
  assign mem[7267] = 10'd6;
  assign mem[7268] = 10'd7;
  assign mem[7269] = 10'd8;
  assign mem[7270] = 10'd2;
  assign mem[7271] = 10'd1;
  assign mem[7272] = 10'd0;
  assign mem[7273] = 10'd1;
  assign mem[7274] = 10'd2;
  assign mem[7275] = 10'd3;
  assign mem[7276] = 10'd4;
  assign mem[7277] = 10'd5;
  assign mem[7278] = 10'd6;
  assign mem[7279] = 10'd7;
  assign mem[7280] = 10'd3;
  assign mem[7281] = 10'd2;
  assign mem[7282] = 10'd1;
  assign mem[7283] = 10'd2;
  assign mem[7284] = 10'd3;
  assign mem[7285] = 10'd4;
  assign mem[7286] = 10'd5;
  assign mem[7287] = 10'd6;
  assign mem[7288] = 10'd7;
  assign mem[7289] = 10'd8;
  assign mem[7290] = 10'd4;
  assign mem[7291] = 10'd3;
  assign mem[7292] = 10'd2;
  assign mem[7293] = 10'd3;
  assign mem[7294] = 10'd4;
  assign mem[7295] = 10'd5;
  assign mem[7296] = 10'd6;
  assign mem[7297] = 10'd7;
  assign mem[7298] = 10'd8;
  assign mem[7299] = 10'd9;
  assign mem[7300] = 10'd10;
  assign mem[7301] = 10'd9;
  assign mem[7302] = 10'd8;
  assign mem[7303] = 10'd7;
  assign mem[7304] = 10'd8;
  assign mem[7305] = 10'd9;
  assign mem[7306] = 10'd10;
  assign mem[7307] = 10'd11;
  assign mem[7308] = 10'd12;
  assign mem[7309] = 10'd13;
  assign mem[7310] = 10'd9;
  assign mem[7311] = 10'd8;
  assign mem[7312] = 10'd7;
  assign mem[7313] = 10'd6;
  assign mem[7314] = 10'd7;
  assign mem[7315] = 10'd8;
  assign mem[7316] = 10'd9;
  assign mem[7317] = 10'd10;
  assign mem[7318] = 10'd11;
  assign mem[7319] = 10'd12;
  assign mem[7320] = 10'd8;
  assign mem[7321] = 10'd7;
  assign mem[7322] = 10'd6;
  assign mem[7323] = 10'd5;
  assign mem[7324] = 10'd6;
  assign mem[7325] = 10'd7;
  assign mem[7326] = 10'd8;
  assign mem[7327] = 10'd9;
  assign mem[7328] = 10'd10;
  assign mem[7329] = 10'd11;
  assign mem[7330] = 10'd7;
  assign mem[7331] = 10'd6;
  assign mem[7332] = 10'd5;
  assign mem[7333] = 10'd4;
  assign mem[7334] = 10'd5;
  assign mem[7335] = 10'd6;
  assign mem[7336] = 10'd7;
  assign mem[7337] = 10'd8;
  assign mem[7338] = 10'd9;
  assign mem[7339] = 10'd10;
  assign mem[7340] = 10'd6;
  assign mem[7341] = 10'd5;
  assign mem[7342] = 10'd4;
  assign mem[7343] = 10'd3;
  assign mem[7344] = 10'd4;
  assign mem[7345] = 10'd5;
  assign mem[7346] = 10'd6;
  assign mem[7347] = 10'd7;
  assign mem[7348] = 10'd8;
  assign mem[7349] = 10'd9;
  assign mem[7350] = 10'd5;
  assign mem[7351] = 10'd4;
  assign mem[7352] = 10'd3;
  assign mem[7353] = 10'd2;
  assign mem[7354] = 10'd3;
  assign mem[7355] = 10'd4;
  assign mem[7356] = 10'd5;
  assign mem[7357] = 10'd6;
  assign mem[7358] = 10'd7;
  assign mem[7359] = 10'd8;
  assign mem[7360] = 10'd4;
  assign mem[7361] = 10'd3;
  assign mem[7362] = 10'd2;
  assign mem[7363] = 10'd1;
  assign mem[7364] = 10'd2;
  assign mem[7365] = 10'd3;
  assign mem[7366] = 10'd4;
  assign mem[7367] = 10'd5;
  assign mem[7368] = 10'd6;
  assign mem[7369] = 10'd7;
  assign mem[7370] = 10'd3;
  assign mem[7371] = 10'd2;
  assign mem[7372] = 10'd1;
  assign mem[7373] = 10'd0;
  assign mem[7374] = 10'd1;
  assign mem[7375] = 10'd2;
  assign mem[7376] = 10'd3;
  assign mem[7377] = 10'd4;
  assign mem[7378] = 10'd5;
  assign mem[7379] = 10'd6;
  assign mem[7380] = 10'd4;
  assign mem[7381] = 10'd3;
  assign mem[7382] = 10'd2;
  assign mem[7383] = 10'd1;
  assign mem[7384] = 10'd2;
  assign mem[7385] = 10'd3;
  assign mem[7386] = 10'd4;
  assign mem[7387] = 10'd5;
  assign mem[7388] = 10'd6;
  assign mem[7389] = 10'd7;
  assign mem[7390] = 10'd5;
  assign mem[7391] = 10'd4;
  assign mem[7392] = 10'd3;
  assign mem[7393] = 10'd2;
  assign mem[7394] = 10'd3;
  assign mem[7395] = 10'd4;
  assign mem[7396] = 10'd5;
  assign mem[7397] = 10'd6;
  assign mem[7398] = 10'd7;
  assign mem[7399] = 10'd8;
  assign mem[7400] = 10'd11;
  assign mem[7401] = 10'd10;
  assign mem[7402] = 10'd9;
  assign mem[7403] = 10'd8;
  assign mem[7404] = 10'd7;
  assign mem[7405] = 10'd8;
  assign mem[7406] = 10'd9;
  assign mem[7407] = 10'd10;
  assign mem[7408] = 10'd11;
  assign mem[7409] = 10'd12;
  assign mem[7410] = 10'd10;
  assign mem[7411] = 10'd9;
  assign mem[7412] = 10'd8;
  assign mem[7413] = 10'd7;
  assign mem[7414] = 10'd6;
  assign mem[7415] = 10'd7;
  assign mem[7416] = 10'd8;
  assign mem[7417] = 10'd9;
  assign mem[7418] = 10'd10;
  assign mem[7419] = 10'd11;
  assign mem[7420] = 10'd9;
  assign mem[7421] = 10'd8;
  assign mem[7422] = 10'd7;
  assign mem[7423] = 10'd6;
  assign mem[7424] = 10'd5;
  assign mem[7425] = 10'd6;
  assign mem[7426] = 10'd7;
  assign mem[7427] = 10'd8;
  assign mem[7428] = 10'd9;
  assign mem[7429] = 10'd10;
  assign mem[7430] = 10'd8;
  assign mem[7431] = 10'd7;
  assign mem[7432] = 10'd6;
  assign mem[7433] = 10'd5;
  assign mem[7434] = 10'd4;
  assign mem[7435] = 10'd5;
  assign mem[7436] = 10'd6;
  assign mem[7437] = 10'd7;
  assign mem[7438] = 10'd8;
  assign mem[7439] = 10'd9;
  assign mem[7440] = 10'd7;
  assign mem[7441] = 10'd6;
  assign mem[7442] = 10'd5;
  assign mem[7443] = 10'd4;
  assign mem[7444] = 10'd3;
  assign mem[7445] = 10'd4;
  assign mem[7446] = 10'd5;
  assign mem[7447] = 10'd6;
  assign mem[7448] = 10'd7;
  assign mem[7449] = 10'd8;
  assign mem[7450] = 10'd6;
  assign mem[7451] = 10'd5;
  assign mem[7452] = 10'd4;
  assign mem[7453] = 10'd3;
  assign mem[7454] = 10'd2;
  assign mem[7455] = 10'd3;
  assign mem[7456] = 10'd4;
  assign mem[7457] = 10'd5;
  assign mem[7458] = 10'd6;
  assign mem[7459] = 10'd7;
  assign mem[7460] = 10'd5;
  assign mem[7461] = 10'd4;
  assign mem[7462] = 10'd3;
  assign mem[7463] = 10'd2;
  assign mem[7464] = 10'd1;
  assign mem[7465] = 10'd2;
  assign mem[7466] = 10'd3;
  assign mem[7467] = 10'd4;
  assign mem[7468] = 10'd5;
  assign mem[7469] = 10'd6;
  assign mem[7470] = 10'd4;
  assign mem[7471] = 10'd3;
  assign mem[7472] = 10'd2;
  assign mem[7473] = 10'd1;
  assign mem[7474] = 10'd0;
  assign mem[7475] = 10'd1;
  assign mem[7476] = 10'd2;
  assign mem[7477] = 10'd3;
  assign mem[7478] = 10'd4;
  assign mem[7479] = 10'd5;
  assign mem[7480] = 10'd5;
  assign mem[7481] = 10'd4;
  assign mem[7482] = 10'd3;
  assign mem[7483] = 10'd2;
  assign mem[7484] = 10'd1;
  assign mem[7485] = 10'd2;
  assign mem[7486] = 10'd3;
  assign mem[7487] = 10'd4;
  assign mem[7488] = 10'd5;
  assign mem[7489] = 10'd6;
  assign mem[7490] = 10'd6;
  assign mem[7491] = 10'd5;
  assign mem[7492] = 10'd4;
  assign mem[7493] = 10'd3;
  assign mem[7494] = 10'd2;
  assign mem[7495] = 10'd3;
  assign mem[7496] = 10'd4;
  assign mem[7497] = 10'd5;
  assign mem[7498] = 10'd6;
  assign mem[7499] = 10'd7;
  assign mem[7500] = 10'd12;
  assign mem[7501] = 10'd11;
  assign mem[7502] = 10'd10;
  assign mem[7503] = 10'd9;
  assign mem[7504] = 10'd8;
  assign mem[7505] = 10'd7;
  assign mem[7506] = 10'd8;
  assign mem[7507] = 10'd9;
  assign mem[7508] = 10'd10;
  assign mem[7509] = 10'd11;
  assign mem[7510] = 10'd11;
  assign mem[7511] = 10'd10;
  assign mem[7512] = 10'd9;
  assign mem[7513] = 10'd8;
  assign mem[7514] = 10'd7;
  assign mem[7515] = 10'd6;
  assign mem[7516] = 10'd7;
  assign mem[7517] = 10'd8;
  assign mem[7518] = 10'd9;
  assign mem[7519] = 10'd10;
  assign mem[7520] = 10'd10;
  assign mem[7521] = 10'd9;
  assign mem[7522] = 10'd8;
  assign mem[7523] = 10'd7;
  assign mem[7524] = 10'd6;
  assign mem[7525] = 10'd5;
  assign mem[7526] = 10'd6;
  assign mem[7527] = 10'd7;
  assign mem[7528] = 10'd8;
  assign mem[7529] = 10'd9;
  assign mem[7530] = 10'd9;
  assign mem[7531] = 10'd8;
  assign mem[7532] = 10'd7;
  assign mem[7533] = 10'd6;
  assign mem[7534] = 10'd5;
  assign mem[7535] = 10'd4;
  assign mem[7536] = 10'd5;
  assign mem[7537] = 10'd6;
  assign mem[7538] = 10'd7;
  assign mem[7539] = 10'd8;
  assign mem[7540] = 10'd8;
  assign mem[7541] = 10'd7;
  assign mem[7542] = 10'd6;
  assign mem[7543] = 10'd5;
  assign mem[7544] = 10'd4;
  assign mem[7545] = 10'd3;
  assign mem[7546] = 10'd4;
  assign mem[7547] = 10'd5;
  assign mem[7548] = 10'd6;
  assign mem[7549] = 10'd7;
  assign mem[7550] = 10'd7;
  assign mem[7551] = 10'd6;
  assign mem[7552] = 10'd5;
  assign mem[7553] = 10'd4;
  assign mem[7554] = 10'd3;
  assign mem[7555] = 10'd2;
  assign mem[7556] = 10'd3;
  assign mem[7557] = 10'd4;
  assign mem[7558] = 10'd5;
  assign mem[7559] = 10'd6;
  assign mem[7560] = 10'd6;
  assign mem[7561] = 10'd5;
  assign mem[7562] = 10'd4;
  assign mem[7563] = 10'd3;
  assign mem[7564] = 10'd2;
  assign mem[7565] = 10'd1;
  assign mem[7566] = 10'd2;
  assign mem[7567] = 10'd3;
  assign mem[7568] = 10'd4;
  assign mem[7569] = 10'd5;
  assign mem[7570] = 10'd5;
  assign mem[7571] = 10'd4;
  assign mem[7572] = 10'd3;
  assign mem[7573] = 10'd2;
  assign mem[7574] = 10'd1;
  assign mem[7575] = 10'd0;
  assign mem[7576] = 10'd1;
  assign mem[7577] = 10'd2;
  assign mem[7578] = 10'd3;
  assign mem[7579] = 10'd4;
  assign mem[7580] = 10'd6;
  assign mem[7581] = 10'd5;
  assign mem[7582] = 10'd4;
  assign mem[7583] = 10'd3;
  assign mem[7584] = 10'd2;
  assign mem[7585] = 10'd1;
  assign mem[7586] = 10'd2;
  assign mem[7587] = 10'd3;
  assign mem[7588] = 10'd4;
  assign mem[7589] = 10'd5;
  assign mem[7590] = 10'd7;
  assign mem[7591] = 10'd6;
  assign mem[7592] = 10'd5;
  assign mem[7593] = 10'd4;
  assign mem[7594] = 10'd3;
  assign mem[7595] = 10'd2;
  assign mem[7596] = 10'd3;
  assign mem[7597] = 10'd4;
  assign mem[7598] = 10'd5;
  assign mem[7599] = 10'd6;
  assign mem[7600] = 10'd13;
  assign mem[7601] = 10'd12;
  assign mem[7602] = 10'd11;
  assign mem[7603] = 10'd10;
  assign mem[7604] = 10'd9;
  assign mem[7605] = 10'd8;
  assign mem[7606] = 10'd7;
  assign mem[7607] = 10'd8;
  assign mem[7608] = 10'd9;
  assign mem[7609] = 10'd10;
  assign mem[7610] = 10'd12;
  assign mem[7611] = 10'd11;
  assign mem[7612] = 10'd10;
  assign mem[7613] = 10'd9;
  assign mem[7614] = 10'd8;
  assign mem[7615] = 10'd7;
  assign mem[7616] = 10'd6;
  assign mem[7617] = 10'd7;
  assign mem[7618] = 10'd8;
  assign mem[7619] = 10'd9;
  assign mem[7620] = 10'd11;
  assign mem[7621] = 10'd10;
  assign mem[7622] = 10'd9;
  assign mem[7623] = 10'd8;
  assign mem[7624] = 10'd7;
  assign mem[7625] = 10'd6;
  assign mem[7626] = 10'd5;
  assign mem[7627] = 10'd6;
  assign mem[7628] = 10'd7;
  assign mem[7629] = 10'd8;
  assign mem[7630] = 10'd10;
  assign mem[7631] = 10'd9;
  assign mem[7632] = 10'd8;
  assign mem[7633] = 10'd7;
  assign mem[7634] = 10'd6;
  assign mem[7635] = 10'd5;
  assign mem[7636] = 10'd4;
  assign mem[7637] = 10'd5;
  assign mem[7638] = 10'd6;
  assign mem[7639] = 10'd7;
  assign mem[7640] = 10'd9;
  assign mem[7641] = 10'd8;
  assign mem[7642] = 10'd7;
  assign mem[7643] = 10'd6;
  assign mem[7644] = 10'd5;
  assign mem[7645] = 10'd4;
  assign mem[7646] = 10'd3;
  assign mem[7647] = 10'd4;
  assign mem[7648] = 10'd5;
  assign mem[7649] = 10'd6;
  assign mem[7650] = 10'd8;
  assign mem[7651] = 10'd7;
  assign mem[7652] = 10'd6;
  assign mem[7653] = 10'd5;
  assign mem[7654] = 10'd4;
  assign mem[7655] = 10'd3;
  assign mem[7656] = 10'd2;
  assign mem[7657] = 10'd3;
  assign mem[7658] = 10'd4;
  assign mem[7659] = 10'd5;
  assign mem[7660] = 10'd7;
  assign mem[7661] = 10'd6;
  assign mem[7662] = 10'd5;
  assign mem[7663] = 10'd4;
  assign mem[7664] = 10'd3;
  assign mem[7665] = 10'd2;
  assign mem[7666] = 10'd1;
  assign mem[7667] = 10'd2;
  assign mem[7668] = 10'd3;
  assign mem[7669] = 10'd4;
  assign mem[7670] = 10'd6;
  assign mem[7671] = 10'd5;
  assign mem[7672] = 10'd4;
  assign mem[7673] = 10'd3;
  assign mem[7674] = 10'd2;
  assign mem[7675] = 10'd1;
  assign mem[7676] = 10'd0;
  assign mem[7677] = 10'd1;
  assign mem[7678] = 10'd2;
  assign mem[7679] = 10'd3;
  assign mem[7680] = 10'd7;
  assign mem[7681] = 10'd6;
  assign mem[7682] = 10'd5;
  assign mem[7683] = 10'd4;
  assign mem[7684] = 10'd3;
  assign mem[7685] = 10'd2;
  assign mem[7686] = 10'd1;
  assign mem[7687] = 10'd2;
  assign mem[7688] = 10'd3;
  assign mem[7689] = 10'd4;
  assign mem[7690] = 10'd8;
  assign mem[7691] = 10'd7;
  assign mem[7692] = 10'd6;
  assign mem[7693] = 10'd5;
  assign mem[7694] = 10'd4;
  assign mem[7695] = 10'd3;
  assign mem[7696] = 10'd2;
  assign mem[7697] = 10'd3;
  assign mem[7698] = 10'd4;
  assign mem[7699] = 10'd5;
  assign mem[7700] = 10'd14;
  assign mem[7701] = 10'd13;
  assign mem[7702] = 10'd12;
  assign mem[7703] = 10'd11;
  assign mem[7704] = 10'd10;
  assign mem[7705] = 10'd9;
  assign mem[7706] = 10'd8;
  assign mem[7707] = 10'd7;
  assign mem[7708] = 10'd8;
  assign mem[7709] = 10'd9;
  assign mem[7710] = 10'd13;
  assign mem[7711] = 10'd12;
  assign mem[7712] = 10'd11;
  assign mem[7713] = 10'd10;
  assign mem[7714] = 10'd9;
  assign mem[7715] = 10'd8;
  assign mem[7716] = 10'd7;
  assign mem[7717] = 10'd6;
  assign mem[7718] = 10'd7;
  assign mem[7719] = 10'd8;
  assign mem[7720] = 10'd12;
  assign mem[7721] = 10'd11;
  assign mem[7722] = 10'd10;
  assign mem[7723] = 10'd9;
  assign mem[7724] = 10'd8;
  assign mem[7725] = 10'd7;
  assign mem[7726] = 10'd6;
  assign mem[7727] = 10'd5;
  assign mem[7728] = 10'd6;
  assign mem[7729] = 10'd7;
  assign mem[7730] = 10'd11;
  assign mem[7731] = 10'd10;
  assign mem[7732] = 10'd9;
  assign mem[7733] = 10'd8;
  assign mem[7734] = 10'd7;
  assign mem[7735] = 10'd6;
  assign mem[7736] = 10'd5;
  assign mem[7737] = 10'd4;
  assign mem[7738] = 10'd5;
  assign mem[7739] = 10'd6;
  assign mem[7740] = 10'd10;
  assign mem[7741] = 10'd9;
  assign mem[7742] = 10'd8;
  assign mem[7743] = 10'd7;
  assign mem[7744] = 10'd6;
  assign mem[7745] = 10'd5;
  assign mem[7746] = 10'd4;
  assign mem[7747] = 10'd3;
  assign mem[7748] = 10'd4;
  assign mem[7749] = 10'd5;
  assign mem[7750] = 10'd9;
  assign mem[7751] = 10'd8;
  assign mem[7752] = 10'd7;
  assign mem[7753] = 10'd6;
  assign mem[7754] = 10'd5;
  assign mem[7755] = 10'd4;
  assign mem[7756] = 10'd3;
  assign mem[7757] = 10'd2;
  assign mem[7758] = 10'd3;
  assign mem[7759] = 10'd4;
  assign mem[7760] = 10'd8;
  assign mem[7761] = 10'd7;
  assign mem[7762] = 10'd6;
  assign mem[7763] = 10'd5;
  assign mem[7764] = 10'd4;
  assign mem[7765] = 10'd3;
  assign mem[7766] = 10'd2;
  assign mem[7767] = 10'd1;
  assign mem[7768] = 10'd2;
  assign mem[7769] = 10'd3;
  assign mem[7770] = 10'd7;
  assign mem[7771] = 10'd6;
  assign mem[7772] = 10'd5;
  assign mem[7773] = 10'd4;
  assign mem[7774] = 10'd3;
  assign mem[7775] = 10'd2;
  assign mem[7776] = 10'd1;
  assign mem[7777] = 10'd0;
  assign mem[7778] = 10'd1;
  assign mem[7779] = 10'd2;
  assign mem[7780] = 10'd8;
  assign mem[7781] = 10'd7;
  assign mem[7782] = 10'd6;
  assign mem[7783] = 10'd5;
  assign mem[7784] = 10'd4;
  assign mem[7785] = 10'd3;
  assign mem[7786] = 10'd2;
  assign mem[7787] = 10'd1;
  assign mem[7788] = 10'd2;
  assign mem[7789] = 10'd3;
  assign mem[7790] = 10'd9;
  assign mem[7791] = 10'd8;
  assign mem[7792] = 10'd7;
  assign mem[7793] = 10'd6;
  assign mem[7794] = 10'd5;
  assign mem[7795] = 10'd4;
  assign mem[7796] = 10'd3;
  assign mem[7797] = 10'd2;
  assign mem[7798] = 10'd3;
  assign mem[7799] = 10'd4;
  assign mem[7800] = 10'd15;
  assign mem[7801] = 10'd14;
  assign mem[7802] = 10'd13;
  assign mem[7803] = 10'd12;
  assign mem[7804] = 10'd11;
  assign mem[7805] = 10'd10;
  assign mem[7806] = 10'd9;
  assign mem[7807] = 10'd8;
  assign mem[7808] = 10'd7;
  assign mem[7809] = 10'd8;
  assign mem[7810] = 10'd14;
  assign mem[7811] = 10'd13;
  assign mem[7812] = 10'd12;
  assign mem[7813] = 10'd11;
  assign mem[7814] = 10'd10;
  assign mem[7815] = 10'd9;
  assign mem[7816] = 10'd8;
  assign mem[7817] = 10'd7;
  assign mem[7818] = 10'd6;
  assign mem[7819] = 10'd7;
  assign mem[7820] = 10'd13;
  assign mem[7821] = 10'd12;
  assign mem[7822] = 10'd11;
  assign mem[7823] = 10'd10;
  assign mem[7824] = 10'd9;
  assign mem[7825] = 10'd8;
  assign mem[7826] = 10'd7;
  assign mem[7827] = 10'd6;
  assign mem[7828] = 10'd5;
  assign mem[7829] = 10'd6;
  assign mem[7830] = 10'd12;
  assign mem[7831] = 10'd11;
  assign mem[7832] = 10'd10;
  assign mem[7833] = 10'd9;
  assign mem[7834] = 10'd8;
  assign mem[7835] = 10'd7;
  assign mem[7836] = 10'd6;
  assign mem[7837] = 10'd5;
  assign mem[7838] = 10'd4;
  assign mem[7839] = 10'd5;
  assign mem[7840] = 10'd11;
  assign mem[7841] = 10'd10;
  assign mem[7842] = 10'd9;
  assign mem[7843] = 10'd8;
  assign mem[7844] = 10'd7;
  assign mem[7845] = 10'd6;
  assign mem[7846] = 10'd5;
  assign mem[7847] = 10'd4;
  assign mem[7848] = 10'd3;
  assign mem[7849] = 10'd4;
  assign mem[7850] = 10'd10;
  assign mem[7851] = 10'd9;
  assign mem[7852] = 10'd8;
  assign mem[7853] = 10'd7;
  assign mem[7854] = 10'd6;
  assign mem[7855] = 10'd5;
  assign mem[7856] = 10'd4;
  assign mem[7857] = 10'd3;
  assign mem[7858] = 10'd2;
  assign mem[7859] = 10'd3;
  assign mem[7860] = 10'd9;
  assign mem[7861] = 10'd8;
  assign mem[7862] = 10'd7;
  assign mem[7863] = 10'd6;
  assign mem[7864] = 10'd5;
  assign mem[7865] = 10'd4;
  assign mem[7866] = 10'd3;
  assign mem[7867] = 10'd2;
  assign mem[7868] = 10'd1;
  assign mem[7869] = 10'd2;
  assign mem[7870] = 10'd8;
  assign mem[7871] = 10'd7;
  assign mem[7872] = 10'd6;
  assign mem[7873] = 10'd5;
  assign mem[7874] = 10'd4;
  assign mem[7875] = 10'd3;
  assign mem[7876] = 10'd2;
  assign mem[7877] = 10'd1;
  assign mem[7878] = 10'd0;
  assign mem[7879] = 10'd1;
  assign mem[7880] = 10'd9;
  assign mem[7881] = 10'd8;
  assign mem[7882] = 10'd7;
  assign mem[7883] = 10'd6;
  assign mem[7884] = 10'd5;
  assign mem[7885] = 10'd4;
  assign mem[7886] = 10'd3;
  assign mem[7887] = 10'd2;
  assign mem[7888] = 10'd1;
  assign mem[7889] = 10'd2;
  assign mem[7890] = 10'd10;
  assign mem[7891] = 10'd9;
  assign mem[7892] = 10'd8;
  assign mem[7893] = 10'd7;
  assign mem[7894] = 10'd6;
  assign mem[7895] = 10'd5;
  assign mem[7896] = 10'd4;
  assign mem[7897] = 10'd3;
  assign mem[7898] = 10'd2;
  assign mem[7899] = 10'd3;
  assign mem[7900] = 10'd16;
  assign mem[7901] = 10'd15;
  assign mem[7902] = 10'd14;
  assign mem[7903] = 10'd13;
  assign mem[7904] = 10'd12;
  assign mem[7905] = 10'd11;
  assign mem[7906] = 10'd10;
  assign mem[7907] = 10'd9;
  assign mem[7908] = 10'd8;
  assign mem[7909] = 10'd7;
  assign mem[7910] = 10'd15;
  assign mem[7911] = 10'd14;
  assign mem[7912] = 10'd13;
  assign mem[7913] = 10'd12;
  assign mem[7914] = 10'd11;
  assign mem[7915] = 10'd10;
  assign mem[7916] = 10'd9;
  assign mem[7917] = 10'd8;
  assign mem[7918] = 10'd7;
  assign mem[7919] = 10'd6;
  assign mem[7920] = 10'd14;
  assign mem[7921] = 10'd13;
  assign mem[7922] = 10'd12;
  assign mem[7923] = 10'd11;
  assign mem[7924] = 10'd10;
  assign mem[7925] = 10'd9;
  assign mem[7926] = 10'd8;
  assign mem[7927] = 10'd7;
  assign mem[7928] = 10'd6;
  assign mem[7929] = 10'd5;
  assign mem[7930] = 10'd13;
  assign mem[7931] = 10'd12;
  assign mem[7932] = 10'd11;
  assign mem[7933] = 10'd10;
  assign mem[7934] = 10'd9;
  assign mem[7935] = 10'd8;
  assign mem[7936] = 10'd7;
  assign mem[7937] = 10'd6;
  assign mem[7938] = 10'd5;
  assign mem[7939] = 10'd4;
  assign mem[7940] = 10'd12;
  assign mem[7941] = 10'd11;
  assign mem[7942] = 10'd10;
  assign mem[7943] = 10'd9;
  assign mem[7944] = 10'd8;
  assign mem[7945] = 10'd7;
  assign mem[7946] = 10'd6;
  assign mem[7947] = 10'd5;
  assign mem[7948] = 10'd4;
  assign mem[7949] = 10'd3;
  assign mem[7950] = 10'd11;
  assign mem[7951] = 10'd10;
  assign mem[7952] = 10'd9;
  assign mem[7953] = 10'd8;
  assign mem[7954] = 10'd7;
  assign mem[7955] = 10'd6;
  assign mem[7956] = 10'd5;
  assign mem[7957] = 10'd4;
  assign mem[7958] = 10'd3;
  assign mem[7959] = 10'd2;
  assign mem[7960] = 10'd10;
  assign mem[7961] = 10'd9;
  assign mem[7962] = 10'd8;
  assign mem[7963] = 10'd7;
  assign mem[7964] = 10'd6;
  assign mem[7965] = 10'd5;
  assign mem[7966] = 10'd4;
  assign mem[7967] = 10'd3;
  assign mem[7968] = 10'd2;
  assign mem[7969] = 10'd1;
  assign mem[7970] = 10'd9;
  assign mem[7971] = 10'd8;
  assign mem[7972] = 10'd7;
  assign mem[7973] = 10'd6;
  assign mem[7974] = 10'd5;
  assign mem[7975] = 10'd4;
  assign mem[7976] = 10'd3;
  assign mem[7977] = 10'd2;
  assign mem[7978] = 10'd1;
  assign mem[7979] = 10'd0;
  assign mem[7980] = 10'd10;
  assign mem[7981] = 10'd9;
  assign mem[7982] = 10'd8;
  assign mem[7983] = 10'd7;
  assign mem[7984] = 10'd6;
  assign mem[7985] = 10'd5;
  assign mem[7986] = 10'd4;
  assign mem[7987] = 10'd3;
  assign mem[7988] = 10'd2;
  assign mem[7989] = 10'd1;
  assign mem[7990] = 10'd11;
  assign mem[7991] = 10'd10;
  assign mem[7992] = 10'd9;
  assign mem[7993] = 10'd8;
  assign mem[7994] = 10'd7;
  assign mem[7995] = 10'd6;
  assign mem[7996] = 10'd5;
  assign mem[7997] = 10'd4;
  assign mem[7998] = 10'd3;
  assign mem[7999] = 10'd2;
  assign mem[8000] = 10'd8;
  assign mem[8001] = 10'd9;
  assign mem[8002] = 10'd10;
  assign mem[8003] = 10'd11;
  assign mem[8004] = 10'd12;
  assign mem[8005] = 10'd13;
  assign mem[8006] = 10'd14;
  assign mem[8007] = 10'd15;
  assign mem[8008] = 10'd16;
  assign mem[8009] = 10'd17;
  assign mem[8010] = 10'd7;
  assign mem[8011] = 10'd8;
  assign mem[8012] = 10'd9;
  assign mem[8013] = 10'd10;
  assign mem[8014] = 10'd11;
  assign mem[8015] = 10'd12;
  assign mem[8016] = 10'd13;
  assign mem[8017] = 10'd14;
  assign mem[8018] = 10'd15;
  assign mem[8019] = 10'd16;
  assign mem[8020] = 10'd6;
  assign mem[8021] = 10'd7;
  assign mem[8022] = 10'd8;
  assign mem[8023] = 10'd9;
  assign mem[8024] = 10'd10;
  assign mem[8025] = 10'd11;
  assign mem[8026] = 10'd12;
  assign mem[8027] = 10'd13;
  assign mem[8028] = 10'd14;
  assign mem[8029] = 10'd15;
  assign mem[8030] = 10'd5;
  assign mem[8031] = 10'd6;
  assign mem[8032] = 10'd7;
  assign mem[8033] = 10'd8;
  assign mem[8034] = 10'd9;
  assign mem[8035] = 10'd10;
  assign mem[8036] = 10'd11;
  assign mem[8037] = 10'd12;
  assign mem[8038] = 10'd13;
  assign mem[8039] = 10'd14;
  assign mem[8040] = 10'd4;
  assign mem[8041] = 10'd5;
  assign mem[8042] = 10'd6;
  assign mem[8043] = 10'd7;
  assign mem[8044] = 10'd8;
  assign mem[8045] = 10'd9;
  assign mem[8046] = 10'd10;
  assign mem[8047] = 10'd11;
  assign mem[8048] = 10'd12;
  assign mem[8049] = 10'd13;
  assign mem[8050] = 10'd3;
  assign mem[8051] = 10'd4;
  assign mem[8052] = 10'd5;
  assign mem[8053] = 10'd6;
  assign mem[8054] = 10'd7;
  assign mem[8055] = 10'd8;
  assign mem[8056] = 10'd9;
  assign mem[8057] = 10'd10;
  assign mem[8058] = 10'd11;
  assign mem[8059] = 10'd12;
  assign mem[8060] = 10'd2;
  assign mem[8061] = 10'd3;
  assign mem[8062] = 10'd4;
  assign mem[8063] = 10'd5;
  assign mem[8064] = 10'd6;
  assign mem[8065] = 10'd7;
  assign mem[8066] = 10'd8;
  assign mem[8067] = 10'd9;
  assign mem[8068] = 10'd10;
  assign mem[8069] = 10'd11;
  assign mem[8070] = 10'd1;
  assign mem[8071] = 10'd2;
  assign mem[8072] = 10'd3;
  assign mem[8073] = 10'd4;
  assign mem[8074] = 10'd5;
  assign mem[8075] = 10'd6;
  assign mem[8076] = 10'd7;
  assign mem[8077] = 10'd8;
  assign mem[8078] = 10'd9;
  assign mem[8079] = 10'd10;
  assign mem[8080] = 10'd0;
  assign mem[8081] = 10'd1;
  assign mem[8082] = 10'd2;
  assign mem[8083] = 10'd3;
  assign mem[8084] = 10'd4;
  assign mem[8085] = 10'd5;
  assign mem[8086] = 10'd6;
  assign mem[8087] = 10'd7;
  assign mem[8088] = 10'd8;
  assign mem[8089] = 10'd9;
  assign mem[8090] = 10'd1;
  assign mem[8091] = 10'd2;
  assign mem[8092] = 10'd3;
  assign mem[8093] = 10'd4;
  assign mem[8094] = 10'd5;
  assign mem[8095] = 10'd6;
  assign mem[8096] = 10'd7;
  assign mem[8097] = 10'd8;
  assign mem[8098] = 10'd9;
  assign mem[8099] = 10'd10;
  assign mem[8100] = 10'd9;
  assign mem[8101] = 10'd8;
  assign mem[8102] = 10'd9;
  assign mem[8103] = 10'd10;
  assign mem[8104] = 10'd11;
  assign mem[8105] = 10'd12;
  assign mem[8106] = 10'd13;
  assign mem[8107] = 10'd14;
  assign mem[8108] = 10'd15;
  assign mem[8109] = 10'd16;
  assign mem[8110] = 10'd8;
  assign mem[8111] = 10'd7;
  assign mem[8112] = 10'd8;
  assign mem[8113] = 10'd9;
  assign mem[8114] = 10'd10;
  assign mem[8115] = 10'd11;
  assign mem[8116] = 10'd12;
  assign mem[8117] = 10'd13;
  assign mem[8118] = 10'd14;
  assign mem[8119] = 10'd15;
  assign mem[8120] = 10'd7;
  assign mem[8121] = 10'd6;
  assign mem[8122] = 10'd7;
  assign mem[8123] = 10'd8;
  assign mem[8124] = 10'd9;
  assign mem[8125] = 10'd10;
  assign mem[8126] = 10'd11;
  assign mem[8127] = 10'd12;
  assign mem[8128] = 10'd13;
  assign mem[8129] = 10'd14;
  assign mem[8130] = 10'd6;
  assign mem[8131] = 10'd5;
  assign mem[8132] = 10'd6;
  assign mem[8133] = 10'd7;
  assign mem[8134] = 10'd8;
  assign mem[8135] = 10'd9;
  assign mem[8136] = 10'd10;
  assign mem[8137] = 10'd11;
  assign mem[8138] = 10'd12;
  assign mem[8139] = 10'd13;
  assign mem[8140] = 10'd5;
  assign mem[8141] = 10'd4;
  assign mem[8142] = 10'd5;
  assign mem[8143] = 10'd6;
  assign mem[8144] = 10'd7;
  assign mem[8145] = 10'd8;
  assign mem[8146] = 10'd9;
  assign mem[8147] = 10'd10;
  assign mem[8148] = 10'd11;
  assign mem[8149] = 10'd12;
  assign mem[8150] = 10'd4;
  assign mem[8151] = 10'd3;
  assign mem[8152] = 10'd4;
  assign mem[8153] = 10'd5;
  assign mem[8154] = 10'd6;
  assign mem[8155] = 10'd7;
  assign mem[8156] = 10'd8;
  assign mem[8157] = 10'd9;
  assign mem[8158] = 10'd10;
  assign mem[8159] = 10'd11;
  assign mem[8160] = 10'd3;
  assign mem[8161] = 10'd2;
  assign mem[8162] = 10'd3;
  assign mem[8163] = 10'd4;
  assign mem[8164] = 10'd5;
  assign mem[8165] = 10'd6;
  assign mem[8166] = 10'd7;
  assign mem[8167] = 10'd8;
  assign mem[8168] = 10'd9;
  assign mem[8169] = 10'd10;
  assign mem[8170] = 10'd2;
  assign mem[8171] = 10'd1;
  assign mem[8172] = 10'd2;
  assign mem[8173] = 10'd3;
  assign mem[8174] = 10'd4;
  assign mem[8175] = 10'd5;
  assign mem[8176] = 10'd6;
  assign mem[8177] = 10'd7;
  assign mem[8178] = 10'd8;
  assign mem[8179] = 10'd9;
  assign mem[8180] = 10'd1;
  assign mem[8181] = 10'd0;
  assign mem[8182] = 10'd1;
  assign mem[8183] = 10'd2;
  assign mem[8184] = 10'd3;
  assign mem[8185] = 10'd4;
  assign mem[8186] = 10'd5;
  assign mem[8187] = 10'd6;
  assign mem[8188] = 10'd7;
  assign mem[8189] = 10'd8;
  assign mem[8190] = 10'd2;
  assign mem[8191] = 10'd1;
  assign mem[8192] = 10'd2;
  assign mem[8193] = 10'd3;
  assign mem[8194] = 10'd4;
  assign mem[8195] = 10'd5;
  assign mem[8196] = 10'd6;
  assign mem[8197] = 10'd7;
  assign mem[8198] = 10'd8;
  assign mem[8199] = 10'd9;
  assign mem[8200] = 10'd10;
  assign mem[8201] = 10'd9;
  assign mem[8202] = 10'd8;
  assign mem[8203] = 10'd9;
  assign mem[8204] = 10'd10;
  assign mem[8205] = 10'd11;
  assign mem[8206] = 10'd12;
  assign mem[8207] = 10'd13;
  assign mem[8208] = 10'd14;
  assign mem[8209] = 10'd15;
  assign mem[8210] = 10'd9;
  assign mem[8211] = 10'd8;
  assign mem[8212] = 10'd7;
  assign mem[8213] = 10'd8;
  assign mem[8214] = 10'd9;
  assign mem[8215] = 10'd10;
  assign mem[8216] = 10'd11;
  assign mem[8217] = 10'd12;
  assign mem[8218] = 10'd13;
  assign mem[8219] = 10'd14;
  assign mem[8220] = 10'd8;
  assign mem[8221] = 10'd7;
  assign mem[8222] = 10'd6;
  assign mem[8223] = 10'd7;
  assign mem[8224] = 10'd8;
  assign mem[8225] = 10'd9;
  assign mem[8226] = 10'd10;
  assign mem[8227] = 10'd11;
  assign mem[8228] = 10'd12;
  assign mem[8229] = 10'd13;
  assign mem[8230] = 10'd7;
  assign mem[8231] = 10'd6;
  assign mem[8232] = 10'd5;
  assign mem[8233] = 10'd6;
  assign mem[8234] = 10'd7;
  assign mem[8235] = 10'd8;
  assign mem[8236] = 10'd9;
  assign mem[8237] = 10'd10;
  assign mem[8238] = 10'd11;
  assign mem[8239] = 10'd12;
  assign mem[8240] = 10'd6;
  assign mem[8241] = 10'd5;
  assign mem[8242] = 10'd4;
  assign mem[8243] = 10'd5;
  assign mem[8244] = 10'd6;
  assign mem[8245] = 10'd7;
  assign mem[8246] = 10'd8;
  assign mem[8247] = 10'd9;
  assign mem[8248] = 10'd10;
  assign mem[8249] = 10'd11;
  assign mem[8250] = 10'd5;
  assign mem[8251] = 10'd4;
  assign mem[8252] = 10'd3;
  assign mem[8253] = 10'd4;
  assign mem[8254] = 10'd5;
  assign mem[8255] = 10'd6;
  assign mem[8256] = 10'd7;
  assign mem[8257] = 10'd8;
  assign mem[8258] = 10'd9;
  assign mem[8259] = 10'd10;
  assign mem[8260] = 10'd4;
  assign mem[8261] = 10'd3;
  assign mem[8262] = 10'd2;
  assign mem[8263] = 10'd3;
  assign mem[8264] = 10'd4;
  assign mem[8265] = 10'd5;
  assign mem[8266] = 10'd6;
  assign mem[8267] = 10'd7;
  assign mem[8268] = 10'd8;
  assign mem[8269] = 10'd9;
  assign mem[8270] = 10'd3;
  assign mem[8271] = 10'd2;
  assign mem[8272] = 10'd1;
  assign mem[8273] = 10'd2;
  assign mem[8274] = 10'd3;
  assign mem[8275] = 10'd4;
  assign mem[8276] = 10'd5;
  assign mem[8277] = 10'd6;
  assign mem[8278] = 10'd7;
  assign mem[8279] = 10'd8;
  assign mem[8280] = 10'd2;
  assign mem[8281] = 10'd1;
  assign mem[8282] = 10'd0;
  assign mem[8283] = 10'd1;
  assign mem[8284] = 10'd2;
  assign mem[8285] = 10'd3;
  assign mem[8286] = 10'd4;
  assign mem[8287] = 10'd5;
  assign mem[8288] = 10'd6;
  assign mem[8289] = 10'd7;
  assign mem[8290] = 10'd3;
  assign mem[8291] = 10'd2;
  assign mem[8292] = 10'd1;
  assign mem[8293] = 10'd2;
  assign mem[8294] = 10'd3;
  assign mem[8295] = 10'd4;
  assign mem[8296] = 10'd5;
  assign mem[8297] = 10'd6;
  assign mem[8298] = 10'd7;
  assign mem[8299] = 10'd8;
  assign mem[8300] = 10'd11;
  assign mem[8301] = 10'd10;
  assign mem[8302] = 10'd9;
  assign mem[8303] = 10'd8;
  assign mem[8304] = 10'd9;
  assign mem[8305] = 10'd10;
  assign mem[8306] = 10'd11;
  assign mem[8307] = 10'd12;
  assign mem[8308] = 10'd13;
  assign mem[8309] = 10'd14;
  assign mem[8310] = 10'd10;
  assign mem[8311] = 10'd9;
  assign mem[8312] = 10'd8;
  assign mem[8313] = 10'd7;
  assign mem[8314] = 10'd8;
  assign mem[8315] = 10'd9;
  assign mem[8316] = 10'd10;
  assign mem[8317] = 10'd11;
  assign mem[8318] = 10'd12;
  assign mem[8319] = 10'd13;
  assign mem[8320] = 10'd9;
  assign mem[8321] = 10'd8;
  assign mem[8322] = 10'd7;
  assign mem[8323] = 10'd6;
  assign mem[8324] = 10'd7;
  assign mem[8325] = 10'd8;
  assign mem[8326] = 10'd9;
  assign mem[8327] = 10'd10;
  assign mem[8328] = 10'd11;
  assign mem[8329] = 10'd12;
  assign mem[8330] = 10'd8;
  assign mem[8331] = 10'd7;
  assign mem[8332] = 10'd6;
  assign mem[8333] = 10'd5;
  assign mem[8334] = 10'd6;
  assign mem[8335] = 10'd7;
  assign mem[8336] = 10'd8;
  assign mem[8337] = 10'd9;
  assign mem[8338] = 10'd10;
  assign mem[8339] = 10'd11;
  assign mem[8340] = 10'd7;
  assign mem[8341] = 10'd6;
  assign mem[8342] = 10'd5;
  assign mem[8343] = 10'd4;
  assign mem[8344] = 10'd5;
  assign mem[8345] = 10'd6;
  assign mem[8346] = 10'd7;
  assign mem[8347] = 10'd8;
  assign mem[8348] = 10'd9;
  assign mem[8349] = 10'd10;
  assign mem[8350] = 10'd6;
  assign mem[8351] = 10'd5;
  assign mem[8352] = 10'd4;
  assign mem[8353] = 10'd3;
  assign mem[8354] = 10'd4;
  assign mem[8355] = 10'd5;
  assign mem[8356] = 10'd6;
  assign mem[8357] = 10'd7;
  assign mem[8358] = 10'd8;
  assign mem[8359] = 10'd9;
  assign mem[8360] = 10'd5;
  assign mem[8361] = 10'd4;
  assign mem[8362] = 10'd3;
  assign mem[8363] = 10'd2;
  assign mem[8364] = 10'd3;
  assign mem[8365] = 10'd4;
  assign mem[8366] = 10'd5;
  assign mem[8367] = 10'd6;
  assign mem[8368] = 10'd7;
  assign mem[8369] = 10'd8;
  assign mem[8370] = 10'd4;
  assign mem[8371] = 10'd3;
  assign mem[8372] = 10'd2;
  assign mem[8373] = 10'd1;
  assign mem[8374] = 10'd2;
  assign mem[8375] = 10'd3;
  assign mem[8376] = 10'd4;
  assign mem[8377] = 10'd5;
  assign mem[8378] = 10'd6;
  assign mem[8379] = 10'd7;
  assign mem[8380] = 10'd3;
  assign mem[8381] = 10'd2;
  assign mem[8382] = 10'd1;
  assign mem[8383] = 10'd0;
  assign mem[8384] = 10'd1;
  assign mem[8385] = 10'd2;
  assign mem[8386] = 10'd3;
  assign mem[8387] = 10'd4;
  assign mem[8388] = 10'd5;
  assign mem[8389] = 10'd6;
  assign mem[8390] = 10'd4;
  assign mem[8391] = 10'd3;
  assign mem[8392] = 10'd2;
  assign mem[8393] = 10'd1;
  assign mem[8394] = 10'd2;
  assign mem[8395] = 10'd3;
  assign mem[8396] = 10'd4;
  assign mem[8397] = 10'd5;
  assign mem[8398] = 10'd6;
  assign mem[8399] = 10'd7;
  assign mem[8400] = 10'd12;
  assign mem[8401] = 10'd11;
  assign mem[8402] = 10'd10;
  assign mem[8403] = 10'd9;
  assign mem[8404] = 10'd8;
  assign mem[8405] = 10'd9;
  assign mem[8406] = 10'd10;
  assign mem[8407] = 10'd11;
  assign mem[8408] = 10'd12;
  assign mem[8409] = 10'd13;
  assign mem[8410] = 10'd11;
  assign mem[8411] = 10'd10;
  assign mem[8412] = 10'd9;
  assign mem[8413] = 10'd8;
  assign mem[8414] = 10'd7;
  assign mem[8415] = 10'd8;
  assign mem[8416] = 10'd9;
  assign mem[8417] = 10'd10;
  assign mem[8418] = 10'd11;
  assign mem[8419] = 10'd12;
  assign mem[8420] = 10'd10;
  assign mem[8421] = 10'd9;
  assign mem[8422] = 10'd8;
  assign mem[8423] = 10'd7;
  assign mem[8424] = 10'd6;
  assign mem[8425] = 10'd7;
  assign mem[8426] = 10'd8;
  assign mem[8427] = 10'd9;
  assign mem[8428] = 10'd10;
  assign mem[8429] = 10'd11;
  assign mem[8430] = 10'd9;
  assign mem[8431] = 10'd8;
  assign mem[8432] = 10'd7;
  assign mem[8433] = 10'd6;
  assign mem[8434] = 10'd5;
  assign mem[8435] = 10'd6;
  assign mem[8436] = 10'd7;
  assign mem[8437] = 10'd8;
  assign mem[8438] = 10'd9;
  assign mem[8439] = 10'd10;
  assign mem[8440] = 10'd8;
  assign mem[8441] = 10'd7;
  assign mem[8442] = 10'd6;
  assign mem[8443] = 10'd5;
  assign mem[8444] = 10'd4;
  assign mem[8445] = 10'd5;
  assign mem[8446] = 10'd6;
  assign mem[8447] = 10'd7;
  assign mem[8448] = 10'd8;
  assign mem[8449] = 10'd9;
  assign mem[8450] = 10'd7;
  assign mem[8451] = 10'd6;
  assign mem[8452] = 10'd5;
  assign mem[8453] = 10'd4;
  assign mem[8454] = 10'd3;
  assign mem[8455] = 10'd4;
  assign mem[8456] = 10'd5;
  assign mem[8457] = 10'd6;
  assign mem[8458] = 10'd7;
  assign mem[8459] = 10'd8;
  assign mem[8460] = 10'd6;
  assign mem[8461] = 10'd5;
  assign mem[8462] = 10'd4;
  assign mem[8463] = 10'd3;
  assign mem[8464] = 10'd2;
  assign mem[8465] = 10'd3;
  assign mem[8466] = 10'd4;
  assign mem[8467] = 10'd5;
  assign mem[8468] = 10'd6;
  assign mem[8469] = 10'd7;
  assign mem[8470] = 10'd5;
  assign mem[8471] = 10'd4;
  assign mem[8472] = 10'd3;
  assign mem[8473] = 10'd2;
  assign mem[8474] = 10'd1;
  assign mem[8475] = 10'd2;
  assign mem[8476] = 10'd3;
  assign mem[8477] = 10'd4;
  assign mem[8478] = 10'd5;
  assign mem[8479] = 10'd6;
  assign mem[8480] = 10'd4;
  assign mem[8481] = 10'd3;
  assign mem[8482] = 10'd2;
  assign mem[8483] = 10'd1;
  assign mem[8484] = 10'd0;
  assign mem[8485] = 10'd1;
  assign mem[8486] = 10'd2;
  assign mem[8487] = 10'd3;
  assign mem[8488] = 10'd4;
  assign mem[8489] = 10'd5;
  assign mem[8490] = 10'd5;
  assign mem[8491] = 10'd4;
  assign mem[8492] = 10'd3;
  assign mem[8493] = 10'd2;
  assign mem[8494] = 10'd1;
  assign mem[8495] = 10'd2;
  assign mem[8496] = 10'd3;
  assign mem[8497] = 10'd4;
  assign mem[8498] = 10'd5;
  assign mem[8499] = 10'd6;
  assign mem[8500] = 10'd13;
  assign mem[8501] = 10'd12;
  assign mem[8502] = 10'd11;
  assign mem[8503] = 10'd10;
  assign mem[8504] = 10'd9;
  assign mem[8505] = 10'd8;
  assign mem[8506] = 10'd9;
  assign mem[8507] = 10'd10;
  assign mem[8508] = 10'd11;
  assign mem[8509] = 10'd12;
  assign mem[8510] = 10'd12;
  assign mem[8511] = 10'd11;
  assign mem[8512] = 10'd10;
  assign mem[8513] = 10'd9;
  assign mem[8514] = 10'd8;
  assign mem[8515] = 10'd7;
  assign mem[8516] = 10'd8;
  assign mem[8517] = 10'd9;
  assign mem[8518] = 10'd10;
  assign mem[8519] = 10'd11;
  assign mem[8520] = 10'd11;
  assign mem[8521] = 10'd10;
  assign mem[8522] = 10'd9;
  assign mem[8523] = 10'd8;
  assign mem[8524] = 10'd7;
  assign mem[8525] = 10'd6;
  assign mem[8526] = 10'd7;
  assign mem[8527] = 10'd8;
  assign mem[8528] = 10'd9;
  assign mem[8529] = 10'd10;
  assign mem[8530] = 10'd10;
  assign mem[8531] = 10'd9;
  assign mem[8532] = 10'd8;
  assign mem[8533] = 10'd7;
  assign mem[8534] = 10'd6;
  assign mem[8535] = 10'd5;
  assign mem[8536] = 10'd6;
  assign mem[8537] = 10'd7;
  assign mem[8538] = 10'd8;
  assign mem[8539] = 10'd9;
  assign mem[8540] = 10'd9;
  assign mem[8541] = 10'd8;
  assign mem[8542] = 10'd7;
  assign mem[8543] = 10'd6;
  assign mem[8544] = 10'd5;
  assign mem[8545] = 10'd4;
  assign mem[8546] = 10'd5;
  assign mem[8547] = 10'd6;
  assign mem[8548] = 10'd7;
  assign mem[8549] = 10'd8;
  assign mem[8550] = 10'd8;
  assign mem[8551] = 10'd7;
  assign mem[8552] = 10'd6;
  assign mem[8553] = 10'd5;
  assign mem[8554] = 10'd4;
  assign mem[8555] = 10'd3;
  assign mem[8556] = 10'd4;
  assign mem[8557] = 10'd5;
  assign mem[8558] = 10'd6;
  assign mem[8559] = 10'd7;
  assign mem[8560] = 10'd7;
  assign mem[8561] = 10'd6;
  assign mem[8562] = 10'd5;
  assign mem[8563] = 10'd4;
  assign mem[8564] = 10'd3;
  assign mem[8565] = 10'd2;
  assign mem[8566] = 10'd3;
  assign mem[8567] = 10'd4;
  assign mem[8568] = 10'd5;
  assign mem[8569] = 10'd6;
  assign mem[8570] = 10'd6;
  assign mem[8571] = 10'd5;
  assign mem[8572] = 10'd4;
  assign mem[8573] = 10'd3;
  assign mem[8574] = 10'd2;
  assign mem[8575] = 10'd1;
  assign mem[8576] = 10'd2;
  assign mem[8577] = 10'd3;
  assign mem[8578] = 10'd4;
  assign mem[8579] = 10'd5;
  assign mem[8580] = 10'd5;
  assign mem[8581] = 10'd4;
  assign mem[8582] = 10'd3;
  assign mem[8583] = 10'd2;
  assign mem[8584] = 10'd1;
  assign mem[8585] = 10'd0;
  assign mem[8586] = 10'd1;
  assign mem[8587] = 10'd2;
  assign mem[8588] = 10'd3;
  assign mem[8589] = 10'd4;
  assign mem[8590] = 10'd6;
  assign mem[8591] = 10'd5;
  assign mem[8592] = 10'd4;
  assign mem[8593] = 10'd3;
  assign mem[8594] = 10'd2;
  assign mem[8595] = 10'd1;
  assign mem[8596] = 10'd2;
  assign mem[8597] = 10'd3;
  assign mem[8598] = 10'd4;
  assign mem[8599] = 10'd5;
  assign mem[8600] = 10'd14;
  assign mem[8601] = 10'd13;
  assign mem[8602] = 10'd12;
  assign mem[8603] = 10'd11;
  assign mem[8604] = 10'd10;
  assign mem[8605] = 10'd9;
  assign mem[8606] = 10'd8;
  assign mem[8607] = 10'd9;
  assign mem[8608] = 10'd10;
  assign mem[8609] = 10'd11;
  assign mem[8610] = 10'd13;
  assign mem[8611] = 10'd12;
  assign mem[8612] = 10'd11;
  assign mem[8613] = 10'd10;
  assign mem[8614] = 10'd9;
  assign mem[8615] = 10'd8;
  assign mem[8616] = 10'd7;
  assign mem[8617] = 10'd8;
  assign mem[8618] = 10'd9;
  assign mem[8619] = 10'd10;
  assign mem[8620] = 10'd12;
  assign mem[8621] = 10'd11;
  assign mem[8622] = 10'd10;
  assign mem[8623] = 10'd9;
  assign mem[8624] = 10'd8;
  assign mem[8625] = 10'd7;
  assign mem[8626] = 10'd6;
  assign mem[8627] = 10'd7;
  assign mem[8628] = 10'd8;
  assign mem[8629] = 10'd9;
  assign mem[8630] = 10'd11;
  assign mem[8631] = 10'd10;
  assign mem[8632] = 10'd9;
  assign mem[8633] = 10'd8;
  assign mem[8634] = 10'd7;
  assign mem[8635] = 10'd6;
  assign mem[8636] = 10'd5;
  assign mem[8637] = 10'd6;
  assign mem[8638] = 10'd7;
  assign mem[8639] = 10'd8;
  assign mem[8640] = 10'd10;
  assign mem[8641] = 10'd9;
  assign mem[8642] = 10'd8;
  assign mem[8643] = 10'd7;
  assign mem[8644] = 10'd6;
  assign mem[8645] = 10'd5;
  assign mem[8646] = 10'd4;
  assign mem[8647] = 10'd5;
  assign mem[8648] = 10'd6;
  assign mem[8649] = 10'd7;
  assign mem[8650] = 10'd9;
  assign mem[8651] = 10'd8;
  assign mem[8652] = 10'd7;
  assign mem[8653] = 10'd6;
  assign mem[8654] = 10'd5;
  assign mem[8655] = 10'd4;
  assign mem[8656] = 10'd3;
  assign mem[8657] = 10'd4;
  assign mem[8658] = 10'd5;
  assign mem[8659] = 10'd6;
  assign mem[8660] = 10'd8;
  assign mem[8661] = 10'd7;
  assign mem[8662] = 10'd6;
  assign mem[8663] = 10'd5;
  assign mem[8664] = 10'd4;
  assign mem[8665] = 10'd3;
  assign mem[8666] = 10'd2;
  assign mem[8667] = 10'd3;
  assign mem[8668] = 10'd4;
  assign mem[8669] = 10'd5;
  assign mem[8670] = 10'd7;
  assign mem[8671] = 10'd6;
  assign mem[8672] = 10'd5;
  assign mem[8673] = 10'd4;
  assign mem[8674] = 10'd3;
  assign mem[8675] = 10'd2;
  assign mem[8676] = 10'd1;
  assign mem[8677] = 10'd2;
  assign mem[8678] = 10'd3;
  assign mem[8679] = 10'd4;
  assign mem[8680] = 10'd6;
  assign mem[8681] = 10'd5;
  assign mem[8682] = 10'd4;
  assign mem[8683] = 10'd3;
  assign mem[8684] = 10'd2;
  assign mem[8685] = 10'd1;
  assign mem[8686] = 10'd0;
  assign mem[8687] = 10'd1;
  assign mem[8688] = 10'd2;
  assign mem[8689] = 10'd3;
  assign mem[8690] = 10'd7;
  assign mem[8691] = 10'd6;
  assign mem[8692] = 10'd5;
  assign mem[8693] = 10'd4;
  assign mem[8694] = 10'd3;
  assign mem[8695] = 10'd2;
  assign mem[8696] = 10'd1;
  assign mem[8697] = 10'd2;
  assign mem[8698] = 10'd3;
  assign mem[8699] = 10'd4;
  assign mem[8700] = 10'd15;
  assign mem[8701] = 10'd14;
  assign mem[8702] = 10'd13;
  assign mem[8703] = 10'd12;
  assign mem[8704] = 10'd11;
  assign mem[8705] = 10'd10;
  assign mem[8706] = 10'd9;
  assign mem[8707] = 10'd8;
  assign mem[8708] = 10'd9;
  assign mem[8709] = 10'd10;
  assign mem[8710] = 10'd14;
  assign mem[8711] = 10'd13;
  assign mem[8712] = 10'd12;
  assign mem[8713] = 10'd11;
  assign mem[8714] = 10'd10;
  assign mem[8715] = 10'd9;
  assign mem[8716] = 10'd8;
  assign mem[8717] = 10'd7;
  assign mem[8718] = 10'd8;
  assign mem[8719] = 10'd9;
  assign mem[8720] = 10'd13;
  assign mem[8721] = 10'd12;
  assign mem[8722] = 10'd11;
  assign mem[8723] = 10'd10;
  assign mem[8724] = 10'd9;
  assign mem[8725] = 10'd8;
  assign mem[8726] = 10'd7;
  assign mem[8727] = 10'd6;
  assign mem[8728] = 10'd7;
  assign mem[8729] = 10'd8;
  assign mem[8730] = 10'd12;
  assign mem[8731] = 10'd11;
  assign mem[8732] = 10'd10;
  assign mem[8733] = 10'd9;
  assign mem[8734] = 10'd8;
  assign mem[8735] = 10'd7;
  assign mem[8736] = 10'd6;
  assign mem[8737] = 10'd5;
  assign mem[8738] = 10'd6;
  assign mem[8739] = 10'd7;
  assign mem[8740] = 10'd11;
  assign mem[8741] = 10'd10;
  assign mem[8742] = 10'd9;
  assign mem[8743] = 10'd8;
  assign mem[8744] = 10'd7;
  assign mem[8745] = 10'd6;
  assign mem[8746] = 10'd5;
  assign mem[8747] = 10'd4;
  assign mem[8748] = 10'd5;
  assign mem[8749] = 10'd6;
  assign mem[8750] = 10'd10;
  assign mem[8751] = 10'd9;
  assign mem[8752] = 10'd8;
  assign mem[8753] = 10'd7;
  assign mem[8754] = 10'd6;
  assign mem[8755] = 10'd5;
  assign mem[8756] = 10'd4;
  assign mem[8757] = 10'd3;
  assign mem[8758] = 10'd4;
  assign mem[8759] = 10'd5;
  assign mem[8760] = 10'd9;
  assign mem[8761] = 10'd8;
  assign mem[8762] = 10'd7;
  assign mem[8763] = 10'd6;
  assign mem[8764] = 10'd5;
  assign mem[8765] = 10'd4;
  assign mem[8766] = 10'd3;
  assign mem[8767] = 10'd2;
  assign mem[8768] = 10'd3;
  assign mem[8769] = 10'd4;
  assign mem[8770] = 10'd8;
  assign mem[8771] = 10'd7;
  assign mem[8772] = 10'd6;
  assign mem[8773] = 10'd5;
  assign mem[8774] = 10'd4;
  assign mem[8775] = 10'd3;
  assign mem[8776] = 10'd2;
  assign mem[8777] = 10'd1;
  assign mem[8778] = 10'd2;
  assign mem[8779] = 10'd3;
  assign mem[8780] = 10'd7;
  assign mem[8781] = 10'd6;
  assign mem[8782] = 10'd5;
  assign mem[8783] = 10'd4;
  assign mem[8784] = 10'd3;
  assign mem[8785] = 10'd2;
  assign mem[8786] = 10'd1;
  assign mem[8787] = 10'd0;
  assign mem[8788] = 10'd1;
  assign mem[8789] = 10'd2;
  assign mem[8790] = 10'd8;
  assign mem[8791] = 10'd7;
  assign mem[8792] = 10'd6;
  assign mem[8793] = 10'd5;
  assign mem[8794] = 10'd4;
  assign mem[8795] = 10'd3;
  assign mem[8796] = 10'd2;
  assign mem[8797] = 10'd1;
  assign mem[8798] = 10'd2;
  assign mem[8799] = 10'd3;
  assign mem[8800] = 10'd16;
  assign mem[8801] = 10'd15;
  assign mem[8802] = 10'd14;
  assign mem[8803] = 10'd13;
  assign mem[8804] = 10'd12;
  assign mem[8805] = 10'd11;
  assign mem[8806] = 10'd10;
  assign mem[8807] = 10'd9;
  assign mem[8808] = 10'd8;
  assign mem[8809] = 10'd9;
  assign mem[8810] = 10'd15;
  assign mem[8811] = 10'd14;
  assign mem[8812] = 10'd13;
  assign mem[8813] = 10'd12;
  assign mem[8814] = 10'd11;
  assign mem[8815] = 10'd10;
  assign mem[8816] = 10'd9;
  assign mem[8817] = 10'd8;
  assign mem[8818] = 10'd7;
  assign mem[8819] = 10'd8;
  assign mem[8820] = 10'd14;
  assign mem[8821] = 10'd13;
  assign mem[8822] = 10'd12;
  assign mem[8823] = 10'd11;
  assign mem[8824] = 10'd10;
  assign mem[8825] = 10'd9;
  assign mem[8826] = 10'd8;
  assign mem[8827] = 10'd7;
  assign mem[8828] = 10'd6;
  assign mem[8829] = 10'd7;
  assign mem[8830] = 10'd13;
  assign mem[8831] = 10'd12;
  assign mem[8832] = 10'd11;
  assign mem[8833] = 10'd10;
  assign mem[8834] = 10'd9;
  assign mem[8835] = 10'd8;
  assign mem[8836] = 10'd7;
  assign mem[8837] = 10'd6;
  assign mem[8838] = 10'd5;
  assign mem[8839] = 10'd6;
  assign mem[8840] = 10'd12;
  assign mem[8841] = 10'd11;
  assign mem[8842] = 10'd10;
  assign mem[8843] = 10'd9;
  assign mem[8844] = 10'd8;
  assign mem[8845] = 10'd7;
  assign mem[8846] = 10'd6;
  assign mem[8847] = 10'd5;
  assign mem[8848] = 10'd4;
  assign mem[8849] = 10'd5;
  assign mem[8850] = 10'd11;
  assign mem[8851] = 10'd10;
  assign mem[8852] = 10'd9;
  assign mem[8853] = 10'd8;
  assign mem[8854] = 10'd7;
  assign mem[8855] = 10'd6;
  assign mem[8856] = 10'd5;
  assign mem[8857] = 10'd4;
  assign mem[8858] = 10'd3;
  assign mem[8859] = 10'd4;
  assign mem[8860] = 10'd10;
  assign mem[8861] = 10'd9;
  assign mem[8862] = 10'd8;
  assign mem[8863] = 10'd7;
  assign mem[8864] = 10'd6;
  assign mem[8865] = 10'd5;
  assign mem[8866] = 10'd4;
  assign mem[8867] = 10'd3;
  assign mem[8868] = 10'd2;
  assign mem[8869] = 10'd3;
  assign mem[8870] = 10'd9;
  assign mem[8871] = 10'd8;
  assign mem[8872] = 10'd7;
  assign mem[8873] = 10'd6;
  assign mem[8874] = 10'd5;
  assign mem[8875] = 10'd4;
  assign mem[8876] = 10'd3;
  assign mem[8877] = 10'd2;
  assign mem[8878] = 10'd1;
  assign mem[8879] = 10'd2;
  assign mem[8880] = 10'd8;
  assign mem[8881] = 10'd7;
  assign mem[8882] = 10'd6;
  assign mem[8883] = 10'd5;
  assign mem[8884] = 10'd4;
  assign mem[8885] = 10'd3;
  assign mem[8886] = 10'd2;
  assign mem[8887] = 10'd1;
  assign mem[8888] = 10'd0;
  assign mem[8889] = 10'd1;
  assign mem[8890] = 10'd9;
  assign mem[8891] = 10'd8;
  assign mem[8892] = 10'd7;
  assign mem[8893] = 10'd6;
  assign mem[8894] = 10'd5;
  assign mem[8895] = 10'd4;
  assign mem[8896] = 10'd3;
  assign mem[8897] = 10'd2;
  assign mem[8898] = 10'd1;
  assign mem[8899] = 10'd2;
  assign mem[8900] = 10'd17;
  assign mem[8901] = 10'd16;
  assign mem[8902] = 10'd15;
  assign mem[8903] = 10'd14;
  assign mem[8904] = 10'd13;
  assign mem[8905] = 10'd12;
  assign mem[8906] = 10'd11;
  assign mem[8907] = 10'd10;
  assign mem[8908] = 10'd9;
  assign mem[8909] = 10'd8;
  assign mem[8910] = 10'd16;
  assign mem[8911] = 10'd15;
  assign mem[8912] = 10'd14;
  assign mem[8913] = 10'd13;
  assign mem[8914] = 10'd12;
  assign mem[8915] = 10'd11;
  assign mem[8916] = 10'd10;
  assign mem[8917] = 10'd9;
  assign mem[8918] = 10'd8;
  assign mem[8919] = 10'd7;
  assign mem[8920] = 10'd15;
  assign mem[8921] = 10'd14;
  assign mem[8922] = 10'd13;
  assign mem[8923] = 10'd12;
  assign mem[8924] = 10'd11;
  assign mem[8925] = 10'd10;
  assign mem[8926] = 10'd9;
  assign mem[8927] = 10'd8;
  assign mem[8928] = 10'd7;
  assign mem[8929] = 10'd6;
  assign mem[8930] = 10'd14;
  assign mem[8931] = 10'd13;
  assign mem[8932] = 10'd12;
  assign mem[8933] = 10'd11;
  assign mem[8934] = 10'd10;
  assign mem[8935] = 10'd9;
  assign mem[8936] = 10'd8;
  assign mem[8937] = 10'd7;
  assign mem[8938] = 10'd6;
  assign mem[8939] = 10'd5;
  assign mem[8940] = 10'd13;
  assign mem[8941] = 10'd12;
  assign mem[8942] = 10'd11;
  assign mem[8943] = 10'd10;
  assign mem[8944] = 10'd9;
  assign mem[8945] = 10'd8;
  assign mem[8946] = 10'd7;
  assign mem[8947] = 10'd6;
  assign mem[8948] = 10'd5;
  assign mem[8949] = 10'd4;
  assign mem[8950] = 10'd12;
  assign mem[8951] = 10'd11;
  assign mem[8952] = 10'd10;
  assign mem[8953] = 10'd9;
  assign mem[8954] = 10'd8;
  assign mem[8955] = 10'd7;
  assign mem[8956] = 10'd6;
  assign mem[8957] = 10'd5;
  assign mem[8958] = 10'd4;
  assign mem[8959] = 10'd3;
  assign mem[8960] = 10'd11;
  assign mem[8961] = 10'd10;
  assign mem[8962] = 10'd9;
  assign mem[8963] = 10'd8;
  assign mem[8964] = 10'd7;
  assign mem[8965] = 10'd6;
  assign mem[8966] = 10'd5;
  assign mem[8967] = 10'd4;
  assign mem[8968] = 10'd3;
  assign mem[8969] = 10'd2;
  assign mem[8970] = 10'd10;
  assign mem[8971] = 10'd9;
  assign mem[8972] = 10'd8;
  assign mem[8973] = 10'd7;
  assign mem[8974] = 10'd6;
  assign mem[8975] = 10'd5;
  assign mem[8976] = 10'd4;
  assign mem[8977] = 10'd3;
  assign mem[8978] = 10'd2;
  assign mem[8979] = 10'd1;
  assign mem[8980] = 10'd9;
  assign mem[8981] = 10'd8;
  assign mem[8982] = 10'd7;
  assign mem[8983] = 10'd6;
  assign mem[8984] = 10'd5;
  assign mem[8985] = 10'd4;
  assign mem[8986] = 10'd3;
  assign mem[8987] = 10'd2;
  assign mem[8988] = 10'd1;
  assign mem[8989] = 10'd0;
  assign mem[8990] = 10'd10;
  assign mem[8991] = 10'd9;
  assign mem[8992] = 10'd8;
  assign mem[8993] = 10'd7;
  assign mem[8994] = 10'd6;
  assign mem[8995] = 10'd5;
  assign mem[8996] = 10'd4;
  assign mem[8997] = 10'd3;
  assign mem[8998] = 10'd2;
  assign mem[8999] = 10'd1;
  assign mem[9000] = 10'd9;
  assign mem[9001] = 10'd10;
  assign mem[9002] = 10'd11;
  assign mem[9003] = 10'd12;
  assign mem[9004] = 10'd13;
  assign mem[9005] = 10'd14;
  assign mem[9006] = 10'd15;
  assign mem[9007] = 10'd16;
  assign mem[9008] = 10'd17;
  assign mem[9009] = 10'd18;
  assign mem[9010] = 10'd8;
  assign mem[9011] = 10'd9;
  assign mem[9012] = 10'd10;
  assign mem[9013] = 10'd11;
  assign mem[9014] = 10'd12;
  assign mem[9015] = 10'd13;
  assign mem[9016] = 10'd14;
  assign mem[9017] = 10'd15;
  assign mem[9018] = 10'd16;
  assign mem[9019] = 10'd17;
  assign mem[9020] = 10'd7;
  assign mem[9021] = 10'd8;
  assign mem[9022] = 10'd9;
  assign mem[9023] = 10'd10;
  assign mem[9024] = 10'd11;
  assign mem[9025] = 10'd12;
  assign mem[9026] = 10'd13;
  assign mem[9027] = 10'd14;
  assign mem[9028] = 10'd15;
  assign mem[9029] = 10'd16;
  assign mem[9030] = 10'd6;
  assign mem[9031] = 10'd7;
  assign mem[9032] = 10'd8;
  assign mem[9033] = 10'd9;
  assign mem[9034] = 10'd10;
  assign mem[9035] = 10'd11;
  assign mem[9036] = 10'd12;
  assign mem[9037] = 10'd13;
  assign mem[9038] = 10'd14;
  assign mem[9039] = 10'd15;
  assign mem[9040] = 10'd5;
  assign mem[9041] = 10'd6;
  assign mem[9042] = 10'd7;
  assign mem[9043] = 10'd8;
  assign mem[9044] = 10'd9;
  assign mem[9045] = 10'd10;
  assign mem[9046] = 10'd11;
  assign mem[9047] = 10'd12;
  assign mem[9048] = 10'd13;
  assign mem[9049] = 10'd14;
  assign mem[9050] = 10'd4;
  assign mem[9051] = 10'd5;
  assign mem[9052] = 10'd6;
  assign mem[9053] = 10'd7;
  assign mem[9054] = 10'd8;
  assign mem[9055] = 10'd9;
  assign mem[9056] = 10'd10;
  assign mem[9057] = 10'd11;
  assign mem[9058] = 10'd12;
  assign mem[9059] = 10'd13;
  assign mem[9060] = 10'd3;
  assign mem[9061] = 10'd4;
  assign mem[9062] = 10'd5;
  assign mem[9063] = 10'd6;
  assign mem[9064] = 10'd7;
  assign mem[9065] = 10'd8;
  assign mem[9066] = 10'd9;
  assign mem[9067] = 10'd10;
  assign mem[9068] = 10'd11;
  assign mem[9069] = 10'd12;
  assign mem[9070] = 10'd2;
  assign mem[9071] = 10'd3;
  assign mem[9072] = 10'd4;
  assign mem[9073] = 10'd5;
  assign mem[9074] = 10'd6;
  assign mem[9075] = 10'd7;
  assign mem[9076] = 10'd8;
  assign mem[9077] = 10'd9;
  assign mem[9078] = 10'd10;
  assign mem[9079] = 10'd11;
  assign mem[9080] = 10'd1;
  assign mem[9081] = 10'd2;
  assign mem[9082] = 10'd3;
  assign mem[9083] = 10'd4;
  assign mem[9084] = 10'd5;
  assign mem[9085] = 10'd6;
  assign mem[9086] = 10'd7;
  assign mem[9087] = 10'd8;
  assign mem[9088] = 10'd9;
  assign mem[9089] = 10'd10;
  assign mem[9090] = 10'd0;
  assign mem[9091] = 10'd1;
  assign mem[9092] = 10'd2;
  assign mem[9093] = 10'd3;
  assign mem[9094] = 10'd4;
  assign mem[9095] = 10'd5;
  assign mem[9096] = 10'd6;
  assign mem[9097] = 10'd7;
  assign mem[9098] = 10'd8;
  assign mem[9099] = 10'd9;
  assign mem[9100] = 10'd10;
  assign mem[9101] = 10'd9;
  assign mem[9102] = 10'd10;
  assign mem[9103] = 10'd11;
  assign mem[9104] = 10'd12;
  assign mem[9105] = 10'd13;
  assign mem[9106] = 10'd14;
  assign mem[9107] = 10'd15;
  assign mem[9108] = 10'd16;
  assign mem[9109] = 10'd17;
  assign mem[9110] = 10'd9;
  assign mem[9111] = 10'd8;
  assign mem[9112] = 10'd9;
  assign mem[9113] = 10'd10;
  assign mem[9114] = 10'd11;
  assign mem[9115] = 10'd12;
  assign mem[9116] = 10'd13;
  assign mem[9117] = 10'd14;
  assign mem[9118] = 10'd15;
  assign mem[9119] = 10'd16;
  assign mem[9120] = 10'd8;
  assign mem[9121] = 10'd7;
  assign mem[9122] = 10'd8;
  assign mem[9123] = 10'd9;
  assign mem[9124] = 10'd10;
  assign mem[9125] = 10'd11;
  assign mem[9126] = 10'd12;
  assign mem[9127] = 10'd13;
  assign mem[9128] = 10'd14;
  assign mem[9129] = 10'd15;
  assign mem[9130] = 10'd7;
  assign mem[9131] = 10'd6;
  assign mem[9132] = 10'd7;
  assign mem[9133] = 10'd8;
  assign mem[9134] = 10'd9;
  assign mem[9135] = 10'd10;
  assign mem[9136] = 10'd11;
  assign mem[9137] = 10'd12;
  assign mem[9138] = 10'd13;
  assign mem[9139] = 10'd14;
  assign mem[9140] = 10'd6;
  assign mem[9141] = 10'd5;
  assign mem[9142] = 10'd6;
  assign mem[9143] = 10'd7;
  assign mem[9144] = 10'd8;
  assign mem[9145] = 10'd9;
  assign mem[9146] = 10'd10;
  assign mem[9147] = 10'd11;
  assign mem[9148] = 10'd12;
  assign mem[9149] = 10'd13;
  assign mem[9150] = 10'd5;
  assign mem[9151] = 10'd4;
  assign mem[9152] = 10'd5;
  assign mem[9153] = 10'd6;
  assign mem[9154] = 10'd7;
  assign mem[9155] = 10'd8;
  assign mem[9156] = 10'd9;
  assign mem[9157] = 10'd10;
  assign mem[9158] = 10'd11;
  assign mem[9159] = 10'd12;
  assign mem[9160] = 10'd4;
  assign mem[9161] = 10'd3;
  assign mem[9162] = 10'd4;
  assign mem[9163] = 10'd5;
  assign mem[9164] = 10'd6;
  assign mem[9165] = 10'd7;
  assign mem[9166] = 10'd8;
  assign mem[9167] = 10'd9;
  assign mem[9168] = 10'd10;
  assign mem[9169] = 10'd11;
  assign mem[9170] = 10'd3;
  assign mem[9171] = 10'd2;
  assign mem[9172] = 10'd3;
  assign mem[9173] = 10'd4;
  assign mem[9174] = 10'd5;
  assign mem[9175] = 10'd6;
  assign mem[9176] = 10'd7;
  assign mem[9177] = 10'd8;
  assign mem[9178] = 10'd9;
  assign mem[9179] = 10'd10;
  assign mem[9180] = 10'd2;
  assign mem[9181] = 10'd1;
  assign mem[9182] = 10'd2;
  assign mem[9183] = 10'd3;
  assign mem[9184] = 10'd4;
  assign mem[9185] = 10'd5;
  assign mem[9186] = 10'd6;
  assign mem[9187] = 10'd7;
  assign mem[9188] = 10'd8;
  assign mem[9189] = 10'd9;
  assign mem[9190] = 10'd1;
  assign mem[9191] = 10'd0;
  assign mem[9192] = 10'd1;
  assign mem[9193] = 10'd2;
  assign mem[9194] = 10'd3;
  assign mem[9195] = 10'd4;
  assign mem[9196] = 10'd5;
  assign mem[9197] = 10'd6;
  assign mem[9198] = 10'd7;
  assign mem[9199] = 10'd8;
  assign mem[9200] = 10'd11;
  assign mem[9201] = 10'd10;
  assign mem[9202] = 10'd9;
  assign mem[9203] = 10'd10;
  assign mem[9204] = 10'd11;
  assign mem[9205] = 10'd12;
  assign mem[9206] = 10'd13;
  assign mem[9207] = 10'd14;
  assign mem[9208] = 10'd15;
  assign mem[9209] = 10'd16;
  assign mem[9210] = 10'd10;
  assign mem[9211] = 10'd9;
  assign mem[9212] = 10'd8;
  assign mem[9213] = 10'd9;
  assign mem[9214] = 10'd10;
  assign mem[9215] = 10'd11;
  assign mem[9216] = 10'd12;
  assign mem[9217] = 10'd13;
  assign mem[9218] = 10'd14;
  assign mem[9219] = 10'd15;
  assign mem[9220] = 10'd9;
  assign mem[9221] = 10'd8;
  assign mem[9222] = 10'd7;
  assign mem[9223] = 10'd8;
  assign mem[9224] = 10'd9;
  assign mem[9225] = 10'd10;
  assign mem[9226] = 10'd11;
  assign mem[9227] = 10'd12;
  assign mem[9228] = 10'd13;
  assign mem[9229] = 10'd14;
  assign mem[9230] = 10'd8;
  assign mem[9231] = 10'd7;
  assign mem[9232] = 10'd6;
  assign mem[9233] = 10'd7;
  assign mem[9234] = 10'd8;
  assign mem[9235] = 10'd9;
  assign mem[9236] = 10'd10;
  assign mem[9237] = 10'd11;
  assign mem[9238] = 10'd12;
  assign mem[9239] = 10'd13;
  assign mem[9240] = 10'd7;
  assign mem[9241] = 10'd6;
  assign mem[9242] = 10'd5;
  assign mem[9243] = 10'd6;
  assign mem[9244] = 10'd7;
  assign mem[9245] = 10'd8;
  assign mem[9246] = 10'd9;
  assign mem[9247] = 10'd10;
  assign mem[9248] = 10'd11;
  assign mem[9249] = 10'd12;
  assign mem[9250] = 10'd6;
  assign mem[9251] = 10'd5;
  assign mem[9252] = 10'd4;
  assign mem[9253] = 10'd5;
  assign mem[9254] = 10'd6;
  assign mem[9255] = 10'd7;
  assign mem[9256] = 10'd8;
  assign mem[9257] = 10'd9;
  assign mem[9258] = 10'd10;
  assign mem[9259] = 10'd11;
  assign mem[9260] = 10'd5;
  assign mem[9261] = 10'd4;
  assign mem[9262] = 10'd3;
  assign mem[9263] = 10'd4;
  assign mem[9264] = 10'd5;
  assign mem[9265] = 10'd6;
  assign mem[9266] = 10'd7;
  assign mem[9267] = 10'd8;
  assign mem[9268] = 10'd9;
  assign mem[9269] = 10'd10;
  assign mem[9270] = 10'd4;
  assign mem[9271] = 10'd3;
  assign mem[9272] = 10'd2;
  assign mem[9273] = 10'd3;
  assign mem[9274] = 10'd4;
  assign mem[9275] = 10'd5;
  assign mem[9276] = 10'd6;
  assign mem[9277] = 10'd7;
  assign mem[9278] = 10'd8;
  assign mem[9279] = 10'd9;
  assign mem[9280] = 10'd3;
  assign mem[9281] = 10'd2;
  assign mem[9282] = 10'd1;
  assign mem[9283] = 10'd2;
  assign mem[9284] = 10'd3;
  assign mem[9285] = 10'd4;
  assign mem[9286] = 10'd5;
  assign mem[9287] = 10'd6;
  assign mem[9288] = 10'd7;
  assign mem[9289] = 10'd8;
  assign mem[9290] = 10'd2;
  assign mem[9291] = 10'd1;
  assign mem[9292] = 10'd0;
  assign mem[9293] = 10'd1;
  assign mem[9294] = 10'd2;
  assign mem[9295] = 10'd3;
  assign mem[9296] = 10'd4;
  assign mem[9297] = 10'd5;
  assign mem[9298] = 10'd6;
  assign mem[9299] = 10'd7;
  assign mem[9300] = 10'd12;
  assign mem[9301] = 10'd11;
  assign mem[9302] = 10'd10;
  assign mem[9303] = 10'd9;
  assign mem[9304] = 10'd10;
  assign mem[9305] = 10'd11;
  assign mem[9306] = 10'd12;
  assign mem[9307] = 10'd13;
  assign mem[9308] = 10'd14;
  assign mem[9309] = 10'd15;
  assign mem[9310] = 10'd11;
  assign mem[9311] = 10'd10;
  assign mem[9312] = 10'd9;
  assign mem[9313] = 10'd8;
  assign mem[9314] = 10'd9;
  assign mem[9315] = 10'd10;
  assign mem[9316] = 10'd11;
  assign mem[9317] = 10'd12;
  assign mem[9318] = 10'd13;
  assign mem[9319] = 10'd14;
  assign mem[9320] = 10'd10;
  assign mem[9321] = 10'd9;
  assign mem[9322] = 10'd8;
  assign mem[9323] = 10'd7;
  assign mem[9324] = 10'd8;
  assign mem[9325] = 10'd9;
  assign mem[9326] = 10'd10;
  assign mem[9327] = 10'd11;
  assign mem[9328] = 10'd12;
  assign mem[9329] = 10'd13;
  assign mem[9330] = 10'd9;
  assign mem[9331] = 10'd8;
  assign mem[9332] = 10'd7;
  assign mem[9333] = 10'd6;
  assign mem[9334] = 10'd7;
  assign mem[9335] = 10'd8;
  assign mem[9336] = 10'd9;
  assign mem[9337] = 10'd10;
  assign mem[9338] = 10'd11;
  assign mem[9339] = 10'd12;
  assign mem[9340] = 10'd8;
  assign mem[9341] = 10'd7;
  assign mem[9342] = 10'd6;
  assign mem[9343] = 10'd5;
  assign mem[9344] = 10'd6;
  assign mem[9345] = 10'd7;
  assign mem[9346] = 10'd8;
  assign mem[9347] = 10'd9;
  assign mem[9348] = 10'd10;
  assign mem[9349] = 10'd11;
  assign mem[9350] = 10'd7;
  assign mem[9351] = 10'd6;
  assign mem[9352] = 10'd5;
  assign mem[9353] = 10'd4;
  assign mem[9354] = 10'd5;
  assign mem[9355] = 10'd6;
  assign mem[9356] = 10'd7;
  assign mem[9357] = 10'd8;
  assign mem[9358] = 10'd9;
  assign mem[9359] = 10'd10;
  assign mem[9360] = 10'd6;
  assign mem[9361] = 10'd5;
  assign mem[9362] = 10'd4;
  assign mem[9363] = 10'd3;
  assign mem[9364] = 10'd4;
  assign mem[9365] = 10'd5;
  assign mem[9366] = 10'd6;
  assign mem[9367] = 10'd7;
  assign mem[9368] = 10'd8;
  assign mem[9369] = 10'd9;
  assign mem[9370] = 10'd5;
  assign mem[9371] = 10'd4;
  assign mem[9372] = 10'd3;
  assign mem[9373] = 10'd2;
  assign mem[9374] = 10'd3;
  assign mem[9375] = 10'd4;
  assign mem[9376] = 10'd5;
  assign mem[9377] = 10'd6;
  assign mem[9378] = 10'd7;
  assign mem[9379] = 10'd8;
  assign mem[9380] = 10'd4;
  assign mem[9381] = 10'd3;
  assign mem[9382] = 10'd2;
  assign mem[9383] = 10'd1;
  assign mem[9384] = 10'd2;
  assign mem[9385] = 10'd3;
  assign mem[9386] = 10'd4;
  assign mem[9387] = 10'd5;
  assign mem[9388] = 10'd6;
  assign mem[9389] = 10'd7;
  assign mem[9390] = 10'd3;
  assign mem[9391] = 10'd2;
  assign mem[9392] = 10'd1;
  assign mem[9393] = 10'd0;
  assign mem[9394] = 10'd1;
  assign mem[9395] = 10'd2;
  assign mem[9396] = 10'd3;
  assign mem[9397] = 10'd4;
  assign mem[9398] = 10'd5;
  assign mem[9399] = 10'd6;
  assign mem[9400] = 10'd13;
  assign mem[9401] = 10'd12;
  assign mem[9402] = 10'd11;
  assign mem[9403] = 10'd10;
  assign mem[9404] = 10'd9;
  assign mem[9405] = 10'd10;
  assign mem[9406] = 10'd11;
  assign mem[9407] = 10'd12;
  assign mem[9408] = 10'd13;
  assign mem[9409] = 10'd14;
  assign mem[9410] = 10'd12;
  assign mem[9411] = 10'd11;
  assign mem[9412] = 10'd10;
  assign mem[9413] = 10'd9;
  assign mem[9414] = 10'd8;
  assign mem[9415] = 10'd9;
  assign mem[9416] = 10'd10;
  assign mem[9417] = 10'd11;
  assign mem[9418] = 10'd12;
  assign mem[9419] = 10'd13;
  assign mem[9420] = 10'd11;
  assign mem[9421] = 10'd10;
  assign mem[9422] = 10'd9;
  assign mem[9423] = 10'd8;
  assign mem[9424] = 10'd7;
  assign mem[9425] = 10'd8;
  assign mem[9426] = 10'd9;
  assign mem[9427] = 10'd10;
  assign mem[9428] = 10'd11;
  assign mem[9429] = 10'd12;
  assign mem[9430] = 10'd10;
  assign mem[9431] = 10'd9;
  assign mem[9432] = 10'd8;
  assign mem[9433] = 10'd7;
  assign mem[9434] = 10'd6;
  assign mem[9435] = 10'd7;
  assign mem[9436] = 10'd8;
  assign mem[9437] = 10'd9;
  assign mem[9438] = 10'd10;
  assign mem[9439] = 10'd11;
  assign mem[9440] = 10'd9;
  assign mem[9441] = 10'd8;
  assign mem[9442] = 10'd7;
  assign mem[9443] = 10'd6;
  assign mem[9444] = 10'd5;
  assign mem[9445] = 10'd6;
  assign mem[9446] = 10'd7;
  assign mem[9447] = 10'd8;
  assign mem[9448] = 10'd9;
  assign mem[9449] = 10'd10;
  assign mem[9450] = 10'd8;
  assign mem[9451] = 10'd7;
  assign mem[9452] = 10'd6;
  assign mem[9453] = 10'd5;
  assign mem[9454] = 10'd4;
  assign mem[9455] = 10'd5;
  assign mem[9456] = 10'd6;
  assign mem[9457] = 10'd7;
  assign mem[9458] = 10'd8;
  assign mem[9459] = 10'd9;
  assign mem[9460] = 10'd7;
  assign mem[9461] = 10'd6;
  assign mem[9462] = 10'd5;
  assign mem[9463] = 10'd4;
  assign mem[9464] = 10'd3;
  assign mem[9465] = 10'd4;
  assign mem[9466] = 10'd5;
  assign mem[9467] = 10'd6;
  assign mem[9468] = 10'd7;
  assign mem[9469] = 10'd8;
  assign mem[9470] = 10'd6;
  assign mem[9471] = 10'd5;
  assign mem[9472] = 10'd4;
  assign mem[9473] = 10'd3;
  assign mem[9474] = 10'd2;
  assign mem[9475] = 10'd3;
  assign mem[9476] = 10'd4;
  assign mem[9477] = 10'd5;
  assign mem[9478] = 10'd6;
  assign mem[9479] = 10'd7;
  assign mem[9480] = 10'd5;
  assign mem[9481] = 10'd4;
  assign mem[9482] = 10'd3;
  assign mem[9483] = 10'd2;
  assign mem[9484] = 10'd1;
  assign mem[9485] = 10'd2;
  assign mem[9486] = 10'd3;
  assign mem[9487] = 10'd4;
  assign mem[9488] = 10'd5;
  assign mem[9489] = 10'd6;
  assign mem[9490] = 10'd4;
  assign mem[9491] = 10'd3;
  assign mem[9492] = 10'd2;
  assign mem[9493] = 10'd1;
  assign mem[9494] = 10'd0;
  assign mem[9495] = 10'd1;
  assign mem[9496] = 10'd2;
  assign mem[9497] = 10'd3;
  assign mem[9498] = 10'd4;
  assign mem[9499] = 10'd5;
  assign mem[9500] = 10'd14;
  assign mem[9501] = 10'd13;
  assign mem[9502] = 10'd12;
  assign mem[9503] = 10'd11;
  assign mem[9504] = 10'd10;
  assign mem[9505] = 10'd9;
  assign mem[9506] = 10'd10;
  assign mem[9507] = 10'd11;
  assign mem[9508] = 10'd12;
  assign mem[9509] = 10'd13;
  assign mem[9510] = 10'd13;
  assign mem[9511] = 10'd12;
  assign mem[9512] = 10'd11;
  assign mem[9513] = 10'd10;
  assign mem[9514] = 10'd9;
  assign mem[9515] = 10'd8;
  assign mem[9516] = 10'd9;
  assign mem[9517] = 10'd10;
  assign mem[9518] = 10'd11;
  assign mem[9519] = 10'd12;
  assign mem[9520] = 10'd12;
  assign mem[9521] = 10'd11;
  assign mem[9522] = 10'd10;
  assign mem[9523] = 10'd9;
  assign mem[9524] = 10'd8;
  assign mem[9525] = 10'd7;
  assign mem[9526] = 10'd8;
  assign mem[9527] = 10'd9;
  assign mem[9528] = 10'd10;
  assign mem[9529] = 10'd11;
  assign mem[9530] = 10'd11;
  assign mem[9531] = 10'd10;
  assign mem[9532] = 10'd9;
  assign mem[9533] = 10'd8;
  assign mem[9534] = 10'd7;
  assign mem[9535] = 10'd6;
  assign mem[9536] = 10'd7;
  assign mem[9537] = 10'd8;
  assign mem[9538] = 10'd9;
  assign mem[9539] = 10'd10;
  assign mem[9540] = 10'd10;
  assign mem[9541] = 10'd9;
  assign mem[9542] = 10'd8;
  assign mem[9543] = 10'd7;
  assign mem[9544] = 10'd6;
  assign mem[9545] = 10'd5;
  assign mem[9546] = 10'd6;
  assign mem[9547] = 10'd7;
  assign mem[9548] = 10'd8;
  assign mem[9549] = 10'd9;
  assign mem[9550] = 10'd9;
  assign mem[9551] = 10'd8;
  assign mem[9552] = 10'd7;
  assign mem[9553] = 10'd6;
  assign mem[9554] = 10'd5;
  assign mem[9555] = 10'd4;
  assign mem[9556] = 10'd5;
  assign mem[9557] = 10'd6;
  assign mem[9558] = 10'd7;
  assign mem[9559] = 10'd8;
  assign mem[9560] = 10'd8;
  assign mem[9561] = 10'd7;
  assign mem[9562] = 10'd6;
  assign mem[9563] = 10'd5;
  assign mem[9564] = 10'd4;
  assign mem[9565] = 10'd3;
  assign mem[9566] = 10'd4;
  assign mem[9567] = 10'd5;
  assign mem[9568] = 10'd6;
  assign mem[9569] = 10'd7;
  assign mem[9570] = 10'd7;
  assign mem[9571] = 10'd6;
  assign mem[9572] = 10'd5;
  assign mem[9573] = 10'd4;
  assign mem[9574] = 10'd3;
  assign mem[9575] = 10'd2;
  assign mem[9576] = 10'd3;
  assign mem[9577] = 10'd4;
  assign mem[9578] = 10'd5;
  assign mem[9579] = 10'd6;
  assign mem[9580] = 10'd6;
  assign mem[9581] = 10'd5;
  assign mem[9582] = 10'd4;
  assign mem[9583] = 10'd3;
  assign mem[9584] = 10'd2;
  assign mem[9585] = 10'd1;
  assign mem[9586] = 10'd2;
  assign mem[9587] = 10'd3;
  assign mem[9588] = 10'd4;
  assign mem[9589] = 10'd5;
  assign mem[9590] = 10'd5;
  assign mem[9591] = 10'd4;
  assign mem[9592] = 10'd3;
  assign mem[9593] = 10'd2;
  assign mem[9594] = 10'd1;
  assign mem[9595] = 10'd0;
  assign mem[9596] = 10'd1;
  assign mem[9597] = 10'd2;
  assign mem[9598] = 10'd3;
  assign mem[9599] = 10'd4;
  assign mem[9600] = 10'd15;
  assign mem[9601] = 10'd14;
  assign mem[9602] = 10'd13;
  assign mem[9603] = 10'd12;
  assign mem[9604] = 10'd11;
  assign mem[9605] = 10'd10;
  assign mem[9606] = 10'd9;
  assign mem[9607] = 10'd10;
  assign mem[9608] = 10'd11;
  assign mem[9609] = 10'd12;
  assign mem[9610] = 10'd14;
  assign mem[9611] = 10'd13;
  assign mem[9612] = 10'd12;
  assign mem[9613] = 10'd11;
  assign mem[9614] = 10'd10;
  assign mem[9615] = 10'd9;
  assign mem[9616] = 10'd8;
  assign mem[9617] = 10'd9;
  assign mem[9618] = 10'd10;
  assign mem[9619] = 10'd11;
  assign mem[9620] = 10'd13;
  assign mem[9621] = 10'd12;
  assign mem[9622] = 10'd11;
  assign mem[9623] = 10'd10;
  assign mem[9624] = 10'd9;
  assign mem[9625] = 10'd8;
  assign mem[9626] = 10'd7;
  assign mem[9627] = 10'd8;
  assign mem[9628] = 10'd9;
  assign mem[9629] = 10'd10;
  assign mem[9630] = 10'd12;
  assign mem[9631] = 10'd11;
  assign mem[9632] = 10'd10;
  assign mem[9633] = 10'd9;
  assign mem[9634] = 10'd8;
  assign mem[9635] = 10'd7;
  assign mem[9636] = 10'd6;
  assign mem[9637] = 10'd7;
  assign mem[9638] = 10'd8;
  assign mem[9639] = 10'd9;
  assign mem[9640] = 10'd11;
  assign mem[9641] = 10'd10;
  assign mem[9642] = 10'd9;
  assign mem[9643] = 10'd8;
  assign mem[9644] = 10'd7;
  assign mem[9645] = 10'd6;
  assign mem[9646] = 10'd5;
  assign mem[9647] = 10'd6;
  assign mem[9648] = 10'd7;
  assign mem[9649] = 10'd8;
  assign mem[9650] = 10'd10;
  assign mem[9651] = 10'd9;
  assign mem[9652] = 10'd8;
  assign mem[9653] = 10'd7;
  assign mem[9654] = 10'd6;
  assign mem[9655] = 10'd5;
  assign mem[9656] = 10'd4;
  assign mem[9657] = 10'd5;
  assign mem[9658] = 10'd6;
  assign mem[9659] = 10'd7;
  assign mem[9660] = 10'd9;
  assign mem[9661] = 10'd8;
  assign mem[9662] = 10'd7;
  assign mem[9663] = 10'd6;
  assign mem[9664] = 10'd5;
  assign mem[9665] = 10'd4;
  assign mem[9666] = 10'd3;
  assign mem[9667] = 10'd4;
  assign mem[9668] = 10'd5;
  assign mem[9669] = 10'd6;
  assign mem[9670] = 10'd8;
  assign mem[9671] = 10'd7;
  assign mem[9672] = 10'd6;
  assign mem[9673] = 10'd5;
  assign mem[9674] = 10'd4;
  assign mem[9675] = 10'd3;
  assign mem[9676] = 10'd2;
  assign mem[9677] = 10'd3;
  assign mem[9678] = 10'd4;
  assign mem[9679] = 10'd5;
  assign mem[9680] = 10'd7;
  assign mem[9681] = 10'd6;
  assign mem[9682] = 10'd5;
  assign mem[9683] = 10'd4;
  assign mem[9684] = 10'd3;
  assign mem[9685] = 10'd2;
  assign mem[9686] = 10'd1;
  assign mem[9687] = 10'd2;
  assign mem[9688] = 10'd3;
  assign mem[9689] = 10'd4;
  assign mem[9690] = 10'd6;
  assign mem[9691] = 10'd5;
  assign mem[9692] = 10'd4;
  assign mem[9693] = 10'd3;
  assign mem[9694] = 10'd2;
  assign mem[9695] = 10'd1;
  assign mem[9696] = 10'd0;
  assign mem[9697] = 10'd1;
  assign mem[9698] = 10'd2;
  assign mem[9699] = 10'd3;
  assign mem[9700] = 10'd16;
  assign mem[9701] = 10'd15;
  assign mem[9702] = 10'd14;
  assign mem[9703] = 10'd13;
  assign mem[9704] = 10'd12;
  assign mem[9705] = 10'd11;
  assign mem[9706] = 10'd10;
  assign mem[9707] = 10'd9;
  assign mem[9708] = 10'd10;
  assign mem[9709] = 10'd11;
  assign mem[9710] = 10'd15;
  assign mem[9711] = 10'd14;
  assign mem[9712] = 10'd13;
  assign mem[9713] = 10'd12;
  assign mem[9714] = 10'd11;
  assign mem[9715] = 10'd10;
  assign mem[9716] = 10'd9;
  assign mem[9717] = 10'd8;
  assign mem[9718] = 10'd9;
  assign mem[9719] = 10'd10;
  assign mem[9720] = 10'd14;
  assign mem[9721] = 10'd13;
  assign mem[9722] = 10'd12;
  assign mem[9723] = 10'd11;
  assign mem[9724] = 10'd10;
  assign mem[9725] = 10'd9;
  assign mem[9726] = 10'd8;
  assign mem[9727] = 10'd7;
  assign mem[9728] = 10'd8;
  assign mem[9729] = 10'd9;
  assign mem[9730] = 10'd13;
  assign mem[9731] = 10'd12;
  assign mem[9732] = 10'd11;
  assign mem[9733] = 10'd10;
  assign mem[9734] = 10'd9;
  assign mem[9735] = 10'd8;
  assign mem[9736] = 10'd7;
  assign mem[9737] = 10'd6;
  assign mem[9738] = 10'd7;
  assign mem[9739] = 10'd8;
  assign mem[9740] = 10'd12;
  assign mem[9741] = 10'd11;
  assign mem[9742] = 10'd10;
  assign mem[9743] = 10'd9;
  assign mem[9744] = 10'd8;
  assign mem[9745] = 10'd7;
  assign mem[9746] = 10'd6;
  assign mem[9747] = 10'd5;
  assign mem[9748] = 10'd6;
  assign mem[9749] = 10'd7;
  assign mem[9750] = 10'd11;
  assign mem[9751] = 10'd10;
  assign mem[9752] = 10'd9;
  assign mem[9753] = 10'd8;
  assign mem[9754] = 10'd7;
  assign mem[9755] = 10'd6;
  assign mem[9756] = 10'd5;
  assign mem[9757] = 10'd4;
  assign mem[9758] = 10'd5;
  assign mem[9759] = 10'd6;
  assign mem[9760] = 10'd10;
  assign mem[9761] = 10'd9;
  assign mem[9762] = 10'd8;
  assign mem[9763] = 10'd7;
  assign mem[9764] = 10'd6;
  assign mem[9765] = 10'd5;
  assign mem[9766] = 10'd4;
  assign mem[9767] = 10'd3;
  assign mem[9768] = 10'd4;
  assign mem[9769] = 10'd5;
  assign mem[9770] = 10'd9;
  assign mem[9771] = 10'd8;
  assign mem[9772] = 10'd7;
  assign mem[9773] = 10'd6;
  assign mem[9774] = 10'd5;
  assign mem[9775] = 10'd4;
  assign mem[9776] = 10'd3;
  assign mem[9777] = 10'd2;
  assign mem[9778] = 10'd3;
  assign mem[9779] = 10'd4;
  assign mem[9780] = 10'd8;
  assign mem[9781] = 10'd7;
  assign mem[9782] = 10'd6;
  assign mem[9783] = 10'd5;
  assign mem[9784] = 10'd4;
  assign mem[9785] = 10'd3;
  assign mem[9786] = 10'd2;
  assign mem[9787] = 10'd1;
  assign mem[9788] = 10'd2;
  assign mem[9789] = 10'd3;
  assign mem[9790] = 10'd7;
  assign mem[9791] = 10'd6;
  assign mem[9792] = 10'd5;
  assign mem[9793] = 10'd4;
  assign mem[9794] = 10'd3;
  assign mem[9795] = 10'd2;
  assign mem[9796] = 10'd1;
  assign mem[9797] = 10'd0;
  assign mem[9798] = 10'd1;
  assign mem[9799] = 10'd2;
  assign mem[9800] = 10'd17;
  assign mem[9801] = 10'd16;
  assign mem[9802] = 10'd15;
  assign mem[9803] = 10'd14;
  assign mem[9804] = 10'd13;
  assign mem[9805] = 10'd12;
  assign mem[9806] = 10'd11;
  assign mem[9807] = 10'd10;
  assign mem[9808] = 10'd9;
  assign mem[9809] = 10'd10;
  assign mem[9810] = 10'd16;
  assign mem[9811] = 10'd15;
  assign mem[9812] = 10'd14;
  assign mem[9813] = 10'd13;
  assign mem[9814] = 10'd12;
  assign mem[9815] = 10'd11;
  assign mem[9816] = 10'd10;
  assign mem[9817] = 10'd9;
  assign mem[9818] = 10'd8;
  assign mem[9819] = 10'd9;
  assign mem[9820] = 10'd15;
  assign mem[9821] = 10'd14;
  assign mem[9822] = 10'd13;
  assign mem[9823] = 10'd12;
  assign mem[9824] = 10'd11;
  assign mem[9825] = 10'd10;
  assign mem[9826] = 10'd9;
  assign mem[9827] = 10'd8;
  assign mem[9828] = 10'd7;
  assign mem[9829] = 10'd8;
  assign mem[9830] = 10'd14;
  assign mem[9831] = 10'd13;
  assign mem[9832] = 10'd12;
  assign mem[9833] = 10'd11;
  assign mem[9834] = 10'd10;
  assign mem[9835] = 10'd9;
  assign mem[9836] = 10'd8;
  assign mem[9837] = 10'd7;
  assign mem[9838] = 10'd6;
  assign mem[9839] = 10'd7;
  assign mem[9840] = 10'd13;
  assign mem[9841] = 10'd12;
  assign mem[9842] = 10'd11;
  assign mem[9843] = 10'd10;
  assign mem[9844] = 10'd9;
  assign mem[9845] = 10'd8;
  assign mem[9846] = 10'd7;
  assign mem[9847] = 10'd6;
  assign mem[9848] = 10'd5;
  assign mem[9849] = 10'd6;
  assign mem[9850] = 10'd12;
  assign mem[9851] = 10'd11;
  assign mem[9852] = 10'd10;
  assign mem[9853] = 10'd9;
  assign mem[9854] = 10'd8;
  assign mem[9855] = 10'd7;
  assign mem[9856] = 10'd6;
  assign mem[9857] = 10'd5;
  assign mem[9858] = 10'd4;
  assign mem[9859] = 10'd5;
  assign mem[9860] = 10'd11;
  assign mem[9861] = 10'd10;
  assign mem[9862] = 10'd9;
  assign mem[9863] = 10'd8;
  assign mem[9864] = 10'd7;
  assign mem[9865] = 10'd6;
  assign mem[9866] = 10'd5;
  assign mem[9867] = 10'd4;
  assign mem[9868] = 10'd3;
  assign mem[9869] = 10'd4;
  assign mem[9870] = 10'd10;
  assign mem[9871] = 10'd9;
  assign mem[9872] = 10'd8;
  assign mem[9873] = 10'd7;
  assign mem[9874] = 10'd6;
  assign mem[9875] = 10'd5;
  assign mem[9876] = 10'd4;
  assign mem[9877] = 10'd3;
  assign mem[9878] = 10'd2;
  assign mem[9879] = 10'd3;
  assign mem[9880] = 10'd9;
  assign mem[9881] = 10'd8;
  assign mem[9882] = 10'd7;
  assign mem[9883] = 10'd6;
  assign mem[9884] = 10'd5;
  assign mem[9885] = 10'd4;
  assign mem[9886] = 10'd3;
  assign mem[9887] = 10'd2;
  assign mem[9888] = 10'd1;
  assign mem[9889] = 10'd2;
  assign mem[9890] = 10'd8;
  assign mem[9891] = 10'd7;
  assign mem[9892] = 10'd6;
  assign mem[9893] = 10'd5;
  assign mem[9894] = 10'd4;
  assign mem[9895] = 10'd3;
  assign mem[9896] = 10'd2;
  assign mem[9897] = 10'd1;
  assign mem[9898] = 10'd0;
  assign mem[9899] = 10'd1;
  assign mem[9900] = 10'd18;
  assign mem[9901] = 10'd17;
  assign mem[9902] = 10'd16;
  assign mem[9903] = 10'd15;
  assign mem[9904] = 10'd14;
  assign mem[9905] = 10'd13;
  assign mem[9906] = 10'd12;
  assign mem[9907] = 10'd11;
  assign mem[9908] = 10'd10;
  assign mem[9909] = 10'd9;
  assign mem[9910] = 10'd17;
  assign mem[9911] = 10'd16;
  assign mem[9912] = 10'd15;
  assign mem[9913] = 10'd14;
  assign mem[9914] = 10'd13;
  assign mem[9915] = 10'd12;
  assign mem[9916] = 10'd11;
  assign mem[9917] = 10'd10;
  assign mem[9918] = 10'd9;
  assign mem[9919] = 10'd8;
  assign mem[9920] = 10'd16;
  assign mem[9921] = 10'd15;
  assign mem[9922] = 10'd14;
  assign mem[9923] = 10'd13;
  assign mem[9924] = 10'd12;
  assign mem[9925] = 10'd11;
  assign mem[9926] = 10'd10;
  assign mem[9927] = 10'd9;
  assign mem[9928] = 10'd8;
  assign mem[9929] = 10'd7;
  assign mem[9930] = 10'd15;
  assign mem[9931] = 10'd14;
  assign mem[9932] = 10'd13;
  assign mem[9933] = 10'd12;
  assign mem[9934] = 10'd11;
  assign mem[9935] = 10'd10;
  assign mem[9936] = 10'd9;
  assign mem[9937] = 10'd8;
  assign mem[9938] = 10'd7;
  assign mem[9939] = 10'd6;
  assign mem[9940] = 10'd14;
  assign mem[9941] = 10'd13;
  assign mem[9942] = 10'd12;
  assign mem[9943] = 10'd11;
  assign mem[9944] = 10'd10;
  assign mem[9945] = 10'd9;
  assign mem[9946] = 10'd8;
  assign mem[9947] = 10'd7;
  assign mem[9948] = 10'd6;
  assign mem[9949] = 10'd5;
  assign mem[9950] = 10'd13;
  assign mem[9951] = 10'd12;
  assign mem[9952] = 10'd11;
  assign mem[9953] = 10'd10;
  assign mem[9954] = 10'd9;
  assign mem[9955] = 10'd8;
  assign mem[9956] = 10'd7;
  assign mem[9957] = 10'd6;
  assign mem[9958] = 10'd5;
  assign mem[9959] = 10'd4;
  assign mem[9960] = 10'd12;
  assign mem[9961] = 10'd11;
  assign mem[9962] = 10'd10;
  assign mem[9963] = 10'd9;
  assign mem[9964] = 10'd8;
  assign mem[9965] = 10'd7;
  assign mem[9966] = 10'd6;
  assign mem[9967] = 10'd5;
  assign mem[9968] = 10'd4;
  assign mem[9969] = 10'd3;
  assign mem[9970] = 10'd11;
  assign mem[9971] = 10'd10;
  assign mem[9972] = 10'd9;
  assign mem[9973] = 10'd8;
  assign mem[9974] = 10'd7;
  assign mem[9975] = 10'd6;
  assign mem[9976] = 10'd5;
  assign mem[9977] = 10'd4;
  assign mem[9978] = 10'd3;
  assign mem[9979] = 10'd2;
  assign mem[9980] = 10'd10;
  assign mem[9981] = 10'd9;
  assign mem[9982] = 10'd8;
  assign mem[9983] = 10'd7;
  assign mem[9984] = 10'd6;
  assign mem[9985] = 10'd5;
  assign mem[9986] = 10'd4;
  assign mem[9987] = 10'd3;
  assign mem[9988] = 10'd2;
  assign mem[9989] = 10'd1;
  assign mem[9990] = 10'd9;
  assign mem[9991] = 10'd8;
  assign mem[9992] = 10'd7;
  assign mem[9993] = 10'd6;
  assign mem[9994] = 10'd5;
  assign mem[9995] = 10'd4;
  assign mem[9996] = 10'd3;
  assign mem[9997] = 10'd2;
  assign mem[9998] = 10'd1;
  assign mem[9999] = 10'd0;

endmodule



module st5_d2_s1_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [7-1:0] ca_in,
  input [7-1:0] cb_in,
  input [28-1:0] cva_in,
  input [4-1:0] cva_v_in,
  input [28-1:0] cvb_in,
  input [4-1:0] cvb_v_in,
  input [40-1:0] dvac_in,
  input [40-1:0] dvbc_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [20-1:0] dvac_out,
  output reg [20-1:0] dvbc_out,
  output reg [40-1:0] dvas_out,
  output reg [40-1:0] dvbs_out
);

  wire [7-1:0] cas;
  wire [7-1:0] cbs;
  wire [28-1:0] opva;
  wire [28-1:0] opvb;
  wire [20-1:0] dvac_t;
  wire [20-1:0] dvbc_t;
  wire [40-1:0] dvas_t;
  wire [40-1:0] dvbs_t;
  assign cas = cb_in;
  assign cbs = ca_in;
  assign dvac_t[9:0] = dvac_in[9:0] + dvac_in[19:10];
  assign dvac_t[19:10] = dvac_in[29:20] + dvac_in[39:30];
  assign dvbc_t[9:0] = dvbc_in[9:0] + dvbc_in[19:10];
  assign dvbc_t[19:10] = dvbc_in[29:20] + dvbc_in[39:30];
  assign opva[6:0] = (cva_in[6:0] == cas)? cbs : cva_in[6:0];
  assign opva[13:7] = (cva_in[13:7] == cas)? cbs : cva_in[13:7];
  assign opva[20:14] = (cva_in[20:14] == cas)? cbs : cva_in[20:14];
  assign opva[27:21] = (cva_in[27:21] == cas)? cbs : cva_in[27:21];
  assign opvb[6:0] = (cvb_in[6:0] == cbs)? cas : cvb_in[6:0];
  assign opvb[13:7] = (cvb_in[13:7] == cbs)? cas : cvb_in[13:7];
  assign opvb[20:14] = (cvb_in[20:14] == cbs)? cas : cvb_in[20:14];
  assign opvb[27:21] = (cvb_in[27:21] == cbs)? cas : cvb_in[27:21];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  distance_rom_10_10
  distance_rom_10_10_das_0
  (
    .opa0(cas),
    .opa1(opva[6:0]),
    .opav(cva_v_in[0]),
    .opb0(cas),
    .opb1(opva[13:7]),
    .opbv(cva_v_in[1]),
    .da(dvas_t[9:0]),
    .db(dvas_t[19:10])
  );


  distance_rom_10_10
  distance_rom_10_10_das_1
  (
    .opa0(cas),
    .opa1(opva[20:14]),
    .opav(cva_v_in[2]),
    .opb0(cas),
    .opb1(opva[27:21]),
    .opbv(cva_v_in[3]),
    .da(dvas_t[29:20]),
    .db(dvas_t[39:30])
  );


  distance_rom_10_10
  distance_rom_10_10_dbs_0
  (
    .opa0(cbs),
    .opa1(opvb[6:0]),
    .opav(cvb_v_in[0]),
    .opb0(cbs),
    .opb1(opvb[13:7]),
    .opbv(cvb_v_in[1]),
    .da(dvbs_t[9:0]),
    .db(dvbs_t[19:10])
  );


  distance_rom_10_10
  distance_rom_10_10_dbs_1
  (
    .opa0(cbs),
    .opa1(opvb[20:14]),
    .opav(cvb_v_in[2]),
    .opb0(cbs),
    .opb1(opvb[27:21]),
    .opbv(cvb_v_in[3]),
    .da(dvbs_t[29:20]),
    .db(dvbs_t[39:30])
  );


  initial begin
    idx_out = 0;
    v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st6_s2_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [20-1:0] dvac_in,
  input [20-1:0] dvbc_in,
  input [40-1:0] dvas_in,
  input [40-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [10-1:0] dvac_out,
  output reg [10-1:0] dvbc_out,
  output reg [20-1:0] dvas_out,
  output reg [20-1:0] dvbs_out
);

  wire [10-1:0] dvac_t;
  wire [10-1:0] dvbc_t;
  wire [20-1:0] dvas_t;
  wire [20-1:0] dvbs_t;
  assign dvac_t = dvac_in[9:0] + dvac_in[19:10];
  assign dvbc_t = dvbc_in[9:0] + dvbc_in[19:10];
  assign dvas_t[9:0] = dvas_in[9:0] + dvas_in[19:10];
  assign dvas_t[19:10] = dvas_in[29:20] + dvas_in[39:30];
  assign dvbs_t[9:0] = dvbs_in[9:0] + dvbs_in[19:10];
  assign dvbs_t[19:10] = dvbs_in[29:20] + dvbs_in[39:30];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dvac_out <= dvac_t;
    dvbc_out <= dvbc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dvac_out = 0;
    dvbc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st7_s3_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [10-1:0] dvac_in,
  input [10-1:0] dvbc_in,
  input [20-1:0] dvas_in,
  input [20-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [10-1:0] dc_out,
  output reg [10-1:0] dvas_out,
  output reg [10-1:0] dvbs_out
);

  wire [10-1:0] dc_t;
  wire [10-1:0] dvas_t;
  wire [10-1:0] dvbs_t;
  assign dc_t = dvac_in + dvbc_in;
  assign dvas_t = dvas_in[9:0] + dvas_in[19:10];
  assign dvbs_t = dvbs_in[9:0] + dvbs_in[19:10];

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dc_out <= dc_t;
    dvas_out <= dvas_t;
    dvbs_out <= dvbs_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dc_out = 0;
    dvas_out = 0;
    dvbs_out = 0;
  end


endmodule



module st8_s4_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [10-1:0] dc_in,
  input [10-1:0] dvas_in,
  input [10-1:0] dvbs_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg [10-1:0] dc_out,
  output reg [10-1:0] ds_out
);

  wire [10-1:0] ds_t;
  assign ds_t = dvas_in + dvbs_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    dc_out <= dc_in;
    ds_out <= ds_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    dc_out = 0;
    ds_out = 0;
  end


endmodule



module st9_cmp_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input [10-1:0] dc_in,
  input [10-1:0] ds_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg sw_out
);

  wire sw_t;
  assign sw_t = ds_in < dc_in;

  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    sw_out <= sw_t;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    sw_out = 0;
  end


endmodule



module st10_reg_6th_100cells
(
  input clk,
  input [3-1:0] idx_in,
  input v_in,
  input sw_in,
  output reg [3-1:0] idx_out,
  output reg v_out,
  output reg sw_out
);


  always @(posedge clk) begin
    idx_out <= idx_in;
    v_out <= v_in;
    sw_out <= sw_in;
  end


  initial begin
    idx_out = 0;
    v_out = 0;
    sw_out = 0;
  end


endmodule

